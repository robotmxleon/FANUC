��  X>�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A3  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ����AIO_CN�V� l� RA�C�LO�MOD�_TYP@FIR��HAL�>#INw_OU�FAC� �gINTERCEmPfBI�IZ@����ALRM_�RECO"  �� ALM�"ENB����&ON�!� M�DG/ 0 $DEBUG1A(�"d�$3AO� ."���!_IF� �P $ENABEL@C#� P dC#5U5K�!MA�B 4�"�
� OG�f �d PCOUP�LE,   $�!PP_D0CES�0�!e81�!"PC�> Q� � �$SOFT�T_�IDq2TOTAL7_EQ� $�0�0�NO�2U SPI_OINDE]�5Xq2�SCREEN_N�AM� e2SI�GN�0e?w;�0P�K_FI0	�$THKY#GPA�NE�4 � DU/MMY1dJD�!RUE4RA!RG1R�� � $TIT1d ��� �Dd��D� �Di@�D5�F6��F7�F8�F9�G0 �G�GPA�E�GhA�E�G�1�G �F�G1�G2��B!SBN_CF��!	 8� !J� ; 
2L A_CM�NT�$FLAsGS]�CHE"�� � ELLSET�UP 
� $�HOME_ PR�<0%�SMACR=O�RREPR�XD0D+�0��R{�T �UTOB U��0 9DE7VIC�CTI�0�A� �013�`B�S�e#VAL�#ISP�_UNI�U`_D�ODf7{iFR_F �0K%D13��1c��C_WAqda�jO�FF_U0N�DEL�hLF0EaA�a7b�??a�`$C?���PA#E�C#sAT�B�d� W_PLv�0CH/ <� PU�P�B
2ds�`�QgdsDUT�P�HAgpSF����WELDH2/�0 =Lc7w7atAING�0$�r�1�@�D2�4%$AS_LKIN;tE�w�t_�~�2UCC_AS
B�FAIL�DSB�"�FAL0�AB<�0�NRDY��P�z$�YN�Wq<��`DE6r��`���p+�����tSTK��0+�;s7�;sNO�p��[�̈́r��U* Ȁ%� 9 � �� ��q`�G�pC�G�+�U�S_FT�0vpF�ǂG�SSF���PAUS���ON\7xǓHOU�ŕ�MI�0�0ƔSECȲ2�ryi �rHE8K0�v8vGAP�+�r	�I� � GTH�F��D_I���T=  �l�����`�s9!̅0����9!G�UN1����q���#MO� �cE' � [M�c�\���REV�B7���!XI� �R o � OD�PN-��dPM��}#�;�/��"8�� F�q�  �#��0DfT p =E RD_E%�Iq�$FSSB�&$�CHKB�pEdeAG� �p�  "
�Ա� Vt:5���3� �a_EDu � G� C2��qS�`x�vl �d$OP�0r�2�a<�_OK��Y�TP_C� <�d8�vU �PLAC�^�}��p� xaCOMM� �rD|ƒ��0�`��KO]B��BIGALwLOW� (K:�w�0VAR��d!�1B P0BL�0S �� ,K|aԚPS�`�0M_O]=՗_�CCG�`N�!� �� ��_ID_��� �0�� B.��1S� ~�CCBD	D�!��I�����@�Ҍ84_ CCWp�` OcOL
��P'�MM
�zn�CHs$MEAdP��d`T�P�!��TR1Q�a�CN���FS3��ir�!/0_�F��( D�!�� C�FfT X0GR�V0��MCqNFLI���0UJ�����!� SWIl�&"D�N�P�d��pM�� � �0EED��!��wPo��`�PJedV
�&$�p�1�``�P��ELBOF� �=��=�p/0����3P�� ��V�Ft���G� �A0WARNM�`ju���wP��𼠤 CORx-�8`FLTRju/TRAT Tlp� �$ACC�rTB�� ��r$ORI�.&��RT�P�pg�
`CHG@I��"3�T{�1�I �r�1K��� �`���"�Q���HD���a�2
BJ{PC���3�4�5�6*�7�8�9�!��COfS_rt����3�V�OLLE�C��"MULTAI�b
2��A
1�� ��0T_�R  4� STY2�R���).��p��o� |A06Kb�Ib$���Pc���U�TO=�cE�EX�T!Y�
B!�Q �2 
l���a0��Rut`9�����  �"�� �Q����qc?�l�~#!|��1Y�M�
�P8$  lT}R�� " Lqࠊ/��P��`AX$JOB׍����&;IGx# d��? %?78��3�p%���9_MOR��$ et��FN�
CNG&AF�TBA���6䱀JC��9��D@r��1CUR.KPa`/E\1��%��?��ttaoA4��XbJ��_R��|rEC�LJ�r�H�LJ��DA���I�����2G����RfT&�C ��bG����HANC6$LG��iqda��N�*�Ya�Cᇁ�0|rf�R'L±�mTX���nSDB�WnSRA�SnSAZ�`�X��$  ' FCYT��e�_F��Pn�Re�M
P�QIkOh ������1��e����Cg���A���MP�a� ��HK�&AE�Up�p�Q�V�9 �'�  ]PI���CSXC��Zq( �xs��s��T�R�C�cPN����MG�IsGH"��aWIDR��$VT�P��9�E�F�PA cI�X�P,aQ�1u�CUS�T��U��)R"TI�T����%nAIOV����P_�L����* \q���OR��$!�q���-��OeP��jЅpIp�Q�u��J8�
��0��~}pPXWORK��=+�$SK0���niDBT)PTRw�_ , �l@Ab��s�R0�ؠD��A:0�_C����=�+`H�PL�q��R�A�"��#�D��r�����BJ�b��9�����DB�Q2��-�r~qPR��ΰ�
�pct��. p�E�S�a��LӉ�/��b���( ��0��b��Pj� 91%��ENE����� 2D�R��RE\���3HPC� � .$L��/�$Ӄ�����INE�׶�q_D����ROS��E0"2q��f0��p��PAZ�tAsbE�TURN����MR�Q2UR@�CRŐE�WMwp��SIGN�A&rlPA��W�`�0$Pf13$P�P� 2j���!q����!��DQ���f������׶GO_AW;0���vp��qa���CS'���CYx42O�1�8�8�*��2��2�N�@�x�CtDۣDEVIѐ� 5 P $�RBֳ��I�P<.�i�I_BY�q��T�A9�HNDG�6�������b�DSBLr3ͳ��CqܢLe7 H� �� ��TOFB̶�FEБg')�h�ۣ�f8��DO�a�� MC9�"�`�s(r�(��H�PWp���rݡSLA4���9IINP!Ѐ� ж�|ۡ�:D *�SPNp�#�lƍ�1��W�I1��J��Eȅq87�qW��NT�V#��V ��SKI�STE^��b��p�L��aJ_�Sjb_>����SAF�k���_�SVBEXCLUT��po�D�pLX ���YH��%q��I_yV9`�bPPLYj���������_ML���L�VRFY_4D��M�IO�`   P�%`�b�Oe��LS�|b��4}�$�����P�u��l�Y�AU NFzf@�����)��#�cD�4dͰ� S��r�AF� �CPX����&`� 3;j��pTA#����  ���SGN��<��<@3�P��c _�t�a���qd��rt��`UN>�����<@rD�p]�T`����%`�����9�p�pI>�=� @��F��\tG@OTS����|�������l��L�EMr�NIC!>2K�GM A��i�DAY�sLOADЩ��D��5���E�F pXI�?j�d��~cO� ���5��_RTRQU�@ �D����0Q�p ��EԠ��� ?�K�%>`� �� MP*Pp��A�"'; 3B�'��VDUS�U�.�CABU�B`��NS9@ID�1W�R$�Q!`V[�Vq_#� ; �DI@�J$C� /$VS�SE�#T�B3C�A�� ���|�3B�AE_l�;VE�P�0SW!�!�@x�3�2� @�`�OH�@3PP <IRwq3BB�p�=�!U����t"BAS��o'~P�Pn%[�d� B	� ����RQDW]%MS�� �%AXC'�;LIFEC���� ��	2�N14B5��34BChd@/Ź�Cq`ʡaN�4q�6��OVՐ�%6HEh�3BSUP$�1��	2D�_�4j�BH1_!C�5š�7Z�:W�:qa�7�S��"BcXZ�Pʁ4AY2HEC��T�pސ�NM����r0P�dD `�L��@HE�VXCSI�Z?6k0��[�Nh�U7FFI�0��C���������6��zrM�SWJEE 8��K�EYIMAG�TM���S�A5��F���r>ЁOCVIE �q'F 	�PLQ�_��?� 	$�&`KD�G� ��ST��!>R|�FT��FTD FT|� FPEMAILb ��aAL��FAUL�SHR�*�;pCO�U_�p��T��U�I�< $�S_�S�#�ITճBUF@kG�kG@�jp`p�0	B�Tk�C��Rws�PSAV(e�R�+B d�$ Cg�p��P/d_���$̰_�Pec �i#OT����P@����jA�gAX�sq:pX�P��\c_G3
L�YN_e!�pJ0D�f�W�r�d"MO*_0T��F��� 2�H��^ЈqK��ey&^��5r$�)�4��qLa���nq�S�cC_ܐ���K씐pu�t��Rp�A�u�XnqDSP�F6nrPC�{IM5c�s�q�nq�U�w{0때0��PIPR�nsN!Djp�sTH��"ûr� yTߑ�sHSDI�v�ABSC_�9@`�V���x�v��c~����NV��G��~�*@�v�P	F!�`d�s0p�a���SC�\��sMER|��nqFBCMP�ӦmpET�⌐M�BFU�0DU�P?�M�B
�CD�yH��`�S�OR_NO�ዑN� �%�i�cg��PS*f�Cjpv�C���a��d��`U OH ����c d������� }�锍��9�D�P�疮A�7�8䙡9�0��1��1�
�1�1$�11�1�>�1K�1X�2f�2T���2
�2�2$�U21�2>�2K�2X��3f�3�3��
�3��3$�31�3>�3�K�3X�4f�BAEX9T�TP <sK��p<6p�p2ǋ��aFDR�QT�PV��b	2p�v�.	2REM�F��B�OVM�s��A��T7ROV��DT3`��MX��IN��Q0��N�IND���
	�<i��`$DG�a{#���4P5�D���R�IV"�=2BGEA-R�qIO�K��;N0p}ة�(���@�0><Z_MCM@	1�_�F|0UR"�R� ,t� a? �P0�?��!?��EG��~Qa��Re�S� � P�a��RIM��P�SETUP2_ T D �STD6���<����pI�C��a�RBACrGU T[ �RTt)Nz�%��+p�IFI�Q!+p��А��PT�{b7qFLUI1T�V � Y�PUR�!�W2�r<qv��PT�� I��$�S���?x#�JQpCO�w`�cVRT� x�$SHO���SASSY��a?58�W���j��A�W�RFU��	15q��25q���*@�X |�NAV�`��3���*@x�R=1��VISIJ�&��SC���E�c�T\�AV��O���B%EX$P�O��I\ ��FMR2b�Y o�X�}p�bpN t�{ߍߟ߶ơP���%_f�G�_��B���M4�Y�k�DGC{LFR%DGDYLD��7�5!6.�04�a�5 1UZ�@�	� T�FS�`2T[� P!��bs�`$GEX_���1�`�Ā\2�3�5��)G��9\��
���P�WeO�&DEBU1G��"��GRR�sp�U�BKU�O1n�� 0PO� �;)' ��' Mb�L�OO�ci!SM� E�7b[���� _E �] �@h��T�ERM�%^�&+PO�RIBq� _�&PS#M_OpL� `�%$����(a�'��UP>Rb� -����]�#0^��G�:0ELTO{Q�$USE��NFIc1G2��!���$4�_$UFR���$j�A1}0=�� OT��7��TAX�p��3N;STCpPATM�d@��2PTHJ�;�Ep4P_bD�H2ARTP`�R5�PPa{RG1REL<�:�aSHFT?�H1�1�8_N�R�8��&% � $�'H@a�q�8B���bSHI@��U�� JaAYLO ��a�a���Y�1��~�J�ERVA� 3H7Cp�2�����E�����RC�~�AScYM.q~�H1WJ[7��E��1Y�>�U2TCp�a�5�Q=��5aP��@��bFORCp�MK �z!:c���'"`&�0w0�a2 H9Ob�fd Ԟ2��,& X�OCA1E!��$OP����V�t ����P��Pd��`RŃ�aOUx��3e��R�5Ie h|�1��e$PWRL�3IM;e�BR_�S�40��� �3H1UD�a�t�QBte7�$HSu�!�`ADDR2�HB}!G�2�a�a�aTc��R��x�f H!�S ���u��u
�u��SEv��Y�HSvH�MN��g
 `�Pr��T�@OL���F�.`A�K�t ACR�O��Q1��ND_C���i��A�d��ROU	P��R_�н�E �Q1�h�s��y���y ���x
��y��y$�h�A��n���AVED��wX��uPt:h $���P_D�H Y�^RrPRM_���!_HTTP_i�Hx�wi (*�OBJ��l�b��$2�LE�3��`���j � (#��L�_
�Tp#��qS�P�c��KRL{i?HITCOU��3!6�L`��Q��U�`��`SS��J�QUERY_FLA�r�HWR�N1x��kpgPINCP	U����O����Œ�!tƑ/tƑ��IwOLNw�l 8!�yRu��$SLL�$INPUT_&Y$;`�P,��M��SLY�x�m���M�I��C��B�!{IO��F_AShn}�$L��Ӈ��8A�b_1���V���@HY1�̡��|�wUOPeo `�� �2��¼���æ�[`P�c;`
�.�æ;�$���QUJa�p � K�NEaG4�v7k��Da��2J7�s��J8��7�I_1����7_LAB�1�P���ɸ��APHI���Q���D�J7Jy8*é_KEY�� �KǐLM�ONx�q <��X�R����X�WATC�H_��C��i�EL�D��y� �er �@Р1V�wFP{�CT�RCz����LG���s� !�$LG�Z�R��Űc�ƈ���FD��I ����\!���ȍ ���� e�Dqf�ce���e����e�� e���@0J_@�ѐ1�ѫ�ژF�A��׷���Cd(��SB����c�ֈ�������I���؅��֍ �����RS=��0  �(t�LN��<t��7���N�	�[�"��U��i��PLr�h�7DAU��EA��h���T���GH�R �
���BOO ru�� C���`ITp����� ��REC��GSCR��#���DQ�<�r�qMARGX~p #�,���dM�>������W+���}䟣JG=M��MNCH�s���FN�K��PR�G��UF��b@��F�WD��HL��STP��V��� ������RS'	HzP����C�dD1R���_��	U ����^���m�������G��@PO�

���Ң�OC/ ��E]X��TUI��I#�\�7h�Bt�B�� ��<@<���e��<@�9N�q�3ANA��A2�x@VAIɰ�tCL�EAR�FDCS_CHI$�!s�O�MO�SI��S�B�IGN��<��é�r��T�t�DEVa�LLQ��J�BU�FF	1vu�j@T6��$��EM��������A�bwu��j@���zq�POS1
�%2�%3�!���
0x �h��x�Q@5�����IDX�TP�~B?bO� ��1"6S�T�R��YmrD1 _w$ES6CS; ���b6u6z��#��_�y L����`Ϩ�����`Na�eE�p�e��#�_ z ���\ࢀ�r�C ��MC\�{ ��h�CLDP�UTRQLI��Ty�8I&DFLGmr&@�QZCb�Di�ZG��LDZEDDZEORGy�]mB �ظq�`��D!s�D/r9C|�| �G�DD(^5DZES�PT8@`���@TVRCLM�C)T�O�O;Y3�d�M����_�}'�$D�EBUGGu��XD'ATA~�=�T�@��UFE��TmqC�sMI6p^�~ de���!RQ`�G�DS3TB�`0 �V;��XAX-B��WlE/XCES�����R)MZ`^����R-DPS��RSq_�����V�_�P�X�xk
oh
��MJPTmā aK`�����aMICb�� � �0�"�]w�RCT �N�S��fR��gA�jL��bC�`Cs��aUS�ED� O� ��C�URPX_T�Q��PS�ҡA� NpTt�ZER�p�pS�`E�B�_FR(P��8q�vZ_�Ѓt��l�A�PT ;MKmă \����46�UB��LIÁ�sREQUIREl�MO�|O�{�Rߣ��ML�0Mlń @��������s)R� WMNDz�S�"�c��Z��^�D��v�IN8���v�RSM��x� �a�1E�D�wQ�L�PST+� �� 4)�LO�`�$R�I% �%EX��AN�G�"�QAODAQlŇ�P$ql��MF���&�9�2� p�5K�W��VSUP�5z�AFEpRIGG�� � �fP�3V�@�S�3v�4I�ΰ%C3 �����������`���Q�'�PETI^�� ���} IN^"� �t�MD�I��) ��)�iQ&�H􀚱�)�DIAͱ*�AN�SWQ�)��!)�D���)wQO\�P_��+ �aU��Vg�\@��Q8aOD�_{P^ዃ �h�3�}P�	}��ڨPڮ2 ��᠍P٨KExF���-�$B��ͦ�0ND2xkRB�*�2_TX�4�XTRA�V���&�LO��_��Ibl�&�R
k��R�������� �MRR}2�U�0 #|����AQ d$C'ALI�PW�G�ȷ�2� RIN��̳<;$RְSW0GT���ABC$�D_Jp<��qϰ�_J31�
+�1SP����ϰ	P+�R�3Qͦ�d�ϰ���J����BQO�]!IM�dRCSKAPGJ�ģ�~���J��dRQ������������_AZR��#�ELxB!��kQOCMP��,Q71n�RT�QN�~�c1���l�01�p�tc~�Z|�SMGA ��bTJG�0SCL<,`�SPH_�dP�����B�ϰӰRT�ER�̳��I-N��AC�"����հE��Ѣ0_N���� ��$1dQ� �db�f%�DI9�tSDH,`tX����� $Vհw���c$��怳A(� �"B�@R������H �$BE�L4�d���_ACCEL�������`S_R��U`�aT71Z#3OqEX+BL[r �@C����s��Sq��h>���>�3[sRO/a_�!��o�u�R�*p���_MG!$D�D�����$FW��P���������D}E��PPABN�RO��EE��!���8@���!~Q�P��� R1q_԰~P�`C� �~Y���Q �1YN�PA��\��@�\aM�Q�����OL�t�INC��������R����QENCS�԰��R����TPpI�N+2I[r����N�TVE� ̳23�_U���" LOWL�H k�8@�@DF�T�P���0��b9C�MOS  �d��`u�WcSPERC�H  ]Otp��  ����ʑCbTʑIאA�FNr��A[r�L <�Ùg��k�C>&�YTRK��(1AY ��Mstan![r}%r#�pT�xa�80MOM����Rtb�@���T��ȷ0�#@�!��DU��\r�S_BCKLSH_C" 5�P~tpd���4�):s��CLALM�A� d`[5�CHK8@�04�GLRTYΐ�����Ar�_@�s_UM�S��6C�S����3 LMTN�_L�@<��4P��7E�=@�;�0�� E��c��S"FD�P	C��Hn� ����5�C7P]����CN_b�NGS�F�SF���VF�1���zA"��E~HCAT�>SH @�㲤��dq�!�}�0\q}�qГ�PA�4�_P�5�#_����u& ����#�T�5JfqB`̋S.OG�G�"TORQU8 f�q�)��`�r��!���R_W�% n$zѓ�d��e��eUI"kI0kI��F�``a��oh����VC��0)�$�c1�n��o���fJRK�l�b�f�, DB��Mң, M�u�_DL��"GR�V!dt��t���aH�_���cA�HzCOSU{V�UxLN�`x{�e t��zy��zyLa�z�|�ja�eZsp��aMY��q�xar#�i{�TH�ET0INK23���?�~�pCBD�C5B~�CذAS��i�`Ldw���w�D�SB�㜕�O�GTS��C�U��t�`S��ˊ�s$DU�0"'��Ȳ��b ����!QʒZC�!NE��\�I�p�3`�0�$b�3�A7�`�i�8GuRxRqLPHUu>�>�S�e���u���u@>��vۓŚ�vb�V��QVw�t���V��V��UVěVқV��V�V��H��$�����QT����HěHқH��UH�H��Os�O���O-���O��O��O�ěOқO��O�O�vF>�d����uŴu��SPBALANC�E��bALE��H_7�SP�ѕv¤v�>�vPFULC�C°+�C³u�1�P�U�TO_�0�UT1T2����2Ng1�� �ī��E�#����!�T/ O9���`IN�SEG��bREV8��bDIFX%*�1��V�1�K O!B�K1$s�'2�P�r1tLCHWAR���y�ABgQ�%$MECHm��{���6AX{!P)D��Y�e�y�� 
���Q��n�ROB�CR"��ՏB �MS�K_���� P ��_6 R����Z$1�B��)4�c�IN���MTCOM_C�`>���  ���~��$NORE�v��S�e�� 4��PGR�R��FLA���$XYZ_D�Av�3 "�DEBUb�� ��S��� ��$TCOD:1 ���"��� $BUFINDX w���MOR�� H�� ��j6�!� �)4Ҹ���A5��0TA � ���"G� �� $SIMU�L�P��������O�BJE���ADJ�US����AY_It�Q�D��OUT�P���� � _FI�=�T
`������7Ж ����� ��DNQ FRI37T5�RO�P� Ea: ��OPWO�`��},��SYSBUP��$SOPy��`1�
U��PRUN,U�PA"�D��҄~�_��-B� 7�A�B��/@��IMAG�:1�&�P��IM�8�INp� RGOVRD,�����P� ����L_`w��QM�2�@RB@�# ?AMC_EDT��� /@NP�M|�.A� MY19-A � �,SL���{ ���OVSL��wSDIZ DEX�C���C/!�V`�N ��Q� �����
#C�@T�'!���_SET�P�� a@�PF"�� 1RI����\#_q�e'~!q!�M@�ѝ��@ ���T�ЪPATUS>� $TRC(�' ��#BTM�'�!I���4-A�#z�� D�E� ��"Y��Eҷ!��  K0�!EXE� �1q2%2�$bN#�U � UP���415 ISXNN��'�A��a�) �P�Gc�q $SU�B�!��{!�!#JM/PWAIPP��5�LO	@������$�RCVFAIL_C'� �1R ������A�@�D��E�pR_{PL#DBTB�Q��B� BWDF~�UM�P
DIG����PTNLP
DeBR�Ly�P�P�pPE�EDZ0�CHADO!W�P��~���E��D|��1DEFSP�� � L���@q_�@���CUNI�H�'�@h1R,02#L ����P�!�BV�� ���P��� ���}N4�KET&R`���.PPYB� h{ ߀SIZE��Ш� ��QS��OR~#FORMATp��ODCO��Q��EM2���T	SUXh ��	�PLIJB� �$n�OMP_SW)IT��E��W��o��c��`/@J@AL_� ��P�@G��`B�oi�C:�D�$}E41�J3Dh�� T{PPDCK�h��}CO_J3���8bvb�;�.o@m���"`C_TAf w� ���PAY�,:��d_1�j2�c`J3���k�ev�c[�TIA4y5y6:�MOM2�)sIs6shIsCs`�B�0AD)s�mv6smvCsPUx�NRNt�u6s�uCr��R��` I$PI5��e��eO��e�� �e���ez������� �������1�ђ�8_%�CHIGc�C �5�D���D�5@ ���ă��A��A�5SA�M�$� �����5MOV��I�L�/�� N�J�>��H��@�`W� �`J�U Z&pF�`H��H�IN��`� �������2��ؘ��؛��GAMM춿!��$GET��D�dT�
��LIB�R^1|BI��$HIB]0_� J�m�EG�bz�At�����LWo� ������٦���b��r@�!aC@EU�:�  dnI_�W T� b�ha~�B�IsT�mv|A�c �$Qh� 1���I} R���D;�c�f1�4e�L�EE��!θ�h����@MSWFLDM.`SCRn87����N��y2�tA��P��UR	�I���p�S_SAVE_DXRg�`3NO�`C�! a2�dg�K��o�q�i| 
��i"�����@��bH���cD���H��@>� e�Q�I㈈~��~Ĉ@e�a��A�a14�M�ߪ � G�YL(�s��~�=�S��[ U��%@����o�����	�.��W��� �p�V��M�#�CL"�q���%�1�y2�PMX�O"� �� $��l$W w�6���aw��du� �du�du�d0@4��PP��S``XPO�c�aZ���P��z� -���OMp��f����������:pCON���4�a_�2� |ba1�g�Iy��6s�� Csg�"z����<zaE�PA �`��>®A �`���P�Q�PM�Q}U� � 8:P�QCOUr�� QT�HT@HO��l HY�S�PES5�kUE�W ]�jPO�T�  b�PPU�e��"UN� ����0O{�� �P��5I�3|BROOGRA�!��24O �ITİ� �INFO}� ��Q�
)����O�I,� (M�SL�EQ�Ts�T�	� S��4� 4�:PENAB�� PTION#�DM��\�D�GCF��U"�J@a��Q�R������QOS�_ED�0� ��s ��KA�_#l�E檠NU>'8(AUT<��;%COPYA�]0(\,�A��Ms�Nf j+^�PRUT�� m"�N�OU bs�R�GADJ}�yRX_���B$P�&�
�&W�(P�(ܰ�&�Cl� �3EX @YC���1RGNS������LGO �@`NYQ_FREQ�r�W�r�r1�T�LA�ĳi1�!Ds�eCR1EX�w!�IF���NA	�%�4_G��DTATg@�4c�MAIL�W��1аg�!Q�1V�D4ELEMΑ� ��@�FEASI�e�4��P�Ѐ)Bep�[F"{�W�I U�i2j�o2 ӳ�B�ABaA`E� ��VA�FBASKb�EW��qU��� |�$��A�GRMS_TR �Ca���C�㸀��A��D �"H0�����	gB 2� ���䬔MV�BLWR�T������BxW�wȴD�OU���N�F2P�R�В�[GRIyD�BARS�#TY��z�Odp}�)��Ч _�4!0�R�TO���� � 9�POR�c\�vbSRV�0)<d4fDI��T�`UahdP1�rgh�rg4pi5pi�6pi7pi8TaNF�(���� $VACLU�CZ�MD)�a>��� �~���c�1W� AN�Y��b�1R( w1W�T�OTAL��qWsP�W_3I�QmtREG#ENkz�rX�H�0w53"vR TR�C���kq_S]��w�p#V �!
$�r��BEC�P�qVҵR 4sV_H��PDAR��p2�S_�Y����6S,�AR�R�2� �"IG�_SEh�p4bE_�� �C_�V�a�U����_lF�{��SLGj����c5���T�Up^pS��DDE�SaUc��. ހTE|��	p�� !�q�0��qJ����=CIL�_M�4`�ѳ�p�T�QR [��@���V���C��P9�HA��M���V1��V1ɛ2�؛2ɛ3؛3ɛ4؛4ɚI��p��J�1��U���9�INf�VIABb�����Dщ�2��U2��3��3��4��!4��}�|R� Sg����D $MC�_Fu "�J�LPh�g��"HsM��I����S ��[���	�KEEP_HNADD�!H��@R�	C$��0h��Q���i�OKG�� �X�i���1�3i�REM��@h�]qb������U�4�eh�HPWD  �H�SBMSK~bCOLLABT��pe�Iq�2DIT�I0���!��� ,�M�FL��|�r�YNT��V�M�C���lp�UP_DLY}���DELA��^q�2�Y2 ADR��Q�SKIP��� �4,`� O��NT^�����P_� ���� �� �����q�Ɋ!�ɉ`�� �`�ʣ`�ʰ`�ʽ`����`��9	1�J2RT)0�ǖX�@Tl3 ��'���#@D����D�N RDCx�� ���R�RV ��n��R�1��o��OTRG�E�yC�ӫRFLGpL��$OTSPC�11UM_��F�2T�H2N�Qa��� �1� ��EFv! 11�� l��0$�t��,�AT���# S�� v6��� ���! OT���H�����
z�2��ʈ�������� y�3������)�;�M�_� 2z�4��̂�����P������q�5�����@#5GYq�6���|����� +�z�7����p/AS  z�8���v����.� Pz�S�q�  Q{�ph,�|���EJ4ҥ�a;��"Nv�#IOC���)I1 '�=�R��W=Eh�� r U���gHt �<P��"$DSB�0�0�BGs��Cg��"� M�/U�P�)D� PEZ�2ǐMDG7&1�"d� D��7DBG_�PP�TSJ1�qPG/QAP��3����S232�%� �����u��ICE�U�BFp�4��ARI9T4�FqOPB4�&�oFLOWc�TRM �Srͱ�P'�CU�0M�JCUXTA�'�INTERFAC�4ڭ�UBpw�SCH3Q� t9��G1̍�6�$��OM$L��A�PI��@�vPAP�� Ti Cc��p���H�C=�EFA�"�@��";��c� H���p]r ���b m���F0Q ��"Ł  2� �S��~r�	� �$N�B��U�/u7SWp_J��BVDSPNVJOG��p�3��_P��BOAN�К���L�.FK�@�_MIRjQ�4��MT~��SAPp���Y��P�DGQS?��P&�GQ<�0�UBRKHaA�Fb��b�� bʃb9R�P�@$�7S�PBSO�CBV��N>eDV�Y{16"�$SV���DE_OPl�FS�PD_OVR4�d���Dyb|SOR�g Np�fF`�ggPOVjUSF�j���c�Q�F�fE�L�UFR�A�jTODLCH��W�OVxd �gPWv��gS�E�K`vPނ�  @;�TI�N��1$OFS2hpC�@e�WD�a+t`�aJa"�Ud`TRA��2�QFDг�QM�B_C:��rBZPB�a��F��r�q�SV@��q��@���ùbG�w6�XAMC�B_b@�Rr-�_M�p'B3��"�_pT$CA]P3�D:bd�HBK�A�Fy�IO %���!��PPA|���������x8��"_rDVC_|0 w3ꀤA2���a�͠�R��3	�Xp���7@�PxaUw3\P�&CAB��"Q��p�h�p�^�O �UX�F?SUBCPU 2tPS��� г�t�@Ѻ���s�t�"��$HW_C���@ї���q ���$U3��d��ATTR�I�@"�tPCYCL���NECAN��SF�LTR_2_FI`2#9T�68�LP�[�CHK��_SCT6�SF_�F_����*�FS1�r�CH�A�щ���rB�RSDz�1+a�C1� �_T�~�:��s@E)MG ��McTϢ���Ϣ��W�DIA�G�ERAILAC4����M��LO.`\�$Tf2�"�X� m�X��$�PR�SP� �^@��C݁�0	QsF�UNC��6ARI	N�;�$i��A��S_GPO d�	���pr�	�#�r�CBL����:�A3�/�6�/�D�A`
�t�:�3�LD@�@l`����OQ������TI����2Q�$CE_RIA4�2AF��P�3��Jp��T2��C�C
��q�OI��vDF_L�~ r�A�@LM�3F}AE0HRDYO�QrpRG��H��a ||�;�MULSE+�p�C��]`�$J�j�J�b�g�kFAN_�ALMLVC��W{RN��HARD`��F0��2$SHADOW%pb0��v����1q�U_&p��A�U֠RԤ(BTO_SBR�$D�[PM���߃�e�MPINF�]p$�x����RE�G!&��DG��p�V��@#fDAL_N�tFL �^�$M@����c�0tpq�p ;$2!$YM2{A�R*3�� ��SEG� 7Sl`"/�A'0�$Te2]c>��`��UAXEQWRO�BNZREDNVWRdE0a_��0cSY	`�i�`��S��WRIE0B��ST� OS)@`�`E�D K���D%�GPB��^q5��.>�OTO��D JpARYNS8��>�W�PFI�P�S$LwINK*�GTHWM�@T_��^qJ�96^b�XYZ�B�
7�OFFfpW50�� s� OBLPղ`�;q@�@�FI=���7@3ddղfT_J�1�B�bd���8^b�0 �.y�f�C� �VDU|rI�9.��TUR��X�ß�Fs�X��0NFL�� pm�<����3y0^btq 1�D %KsPM��Te3Ƒ��p������|CORQ2�@[Q��֑���PO���N��m%�CYQ��$OVE�!M2MU@o!� �%	�%�&kA�'o��'��$AN�Z�! ��N1�!�P� &��!�%��!�',5	�,5�#[QE)RxQ�	��E-0�p$��j4A1���`-�D{�x�{�AX;s �B{�>���Y�5]��9 ���9���:( �:� �:@� �:_�:��:1� �6;��9;��9;��9;� �9;�I;�I;�,I;��<I;�LIiA]IDEBU�$���U�Q{r{AB{�y��a�#9Vn�� 
(R� �PU֑\W]a\W��\W (\W�\W�\W_\W����k��Y�LA�B�N%��GR�Og�N��W�B_ ;�Q6���c� J�f9apO%5e8�AfAND ���_4X��b18�~g  W����h=��hZ�� �NT��/s�`VEL�A��$�ay��f�SE�RVE�`�� $�� �Aq!pPOmr�p2 	q��`�1��  ]$&rTRQp�
%sd��/p�3w��2�Du���v�_ � l8˰�q�ERR�2�I��`�$�qTOQ�$� Lm��4��v-�eGu%m��  %s��.q� , qHubp��1RA�q 2'� d	����u;p7 ���$� @�4о2 $tOCl�-���  �{CO�UNT��!��SFZN_CFG.qG� 4됺�`�T� �'�Sɐ���r�y�^�� �MPM㠀���H��#�!���F!A��	5���X��� ���q
�x�tt���9Po��`HEL��~��� 5��B�_BAS��RSR��ɰ��S���r��1�wr�2��3��4���5��6��7��8�we�ROO=��p^ f� NL	�qABs�s�s�ACK9VIN27�T����$U�r�ԡ%�_PU{��Ї�OU=�P��R��v�ՠ��6TPFWD�_KAR�q��pR�EtQ�PT ���QUE��-�� z����I��<SR�� ���`��SEMXQ�fQ�m�A܁STY4�SO�.�DI@���ࡩ7�_TM��M�ANRQq�� EN�D$$KEYSWITCH����S���HEzBEATmM �PE?�LE�r(�!`ɸU��F����SX�DO_HOM���O��(�EFf0PAR�������A�C��O]шp�qOV_Mx@���IOCMl��d!��Q�HK�� D}�粀	U�ޢM7𲤵 m�FORC��WAR�M��bS�OM@� G� @T=�U��UPX�1��2��3��}4b�� �S<��O��L����r��U�NLO^��3�E�D� F�NPX_;AS�� 0���|�� �$SIZ���$VA?`�uMU/LTIP�S����A��� � A$m�T��� g�S���'�C�p��FRIF��27�SȠ��ķ�N=Ft�ODBU��``����u`�Ss�n�� xzpSI�r�TE�]"�SGLO�Tf�&��h�c<��P�STMT���P+���BW� Q�S�HOW��0�SV�\0_GĂ� _$�PC`8�\3�1FBZ��P��SP�A?����EpVD��Â��� �|qA00 �d���#���#��#�T�#�5!�6!�7!�U8!�9!�A!�B!�@��#��Q$���#�F!��\@��-�1:�1G�1�T�1a�1n�1{�1���1��1��1��1���1��1��1��2� �2-�2:�2G�2*T�2a�2n�2{�^T���2��2��2��2��2��2����P-�c �G�3T�3a�U3n�3{�3��3��U3��3��3��3��U3��3��4�4-�U4:�4G�4T�4a�U4n�4{�4��4��U4��4��4��4��U4��4��5�5-�U5:�5G�5T�5a�U5n�5{�5��5��U5��5��5��5��U5��5��6�6-�U6:�6G�6T�6a�U6n�6{�6��6��U6��6��6��6��U6��6��7�7-�U7:�7G�7T�7a�U7n�7{�7��7��U7��7��7��7��e7��7���rVPǰ=U,r� 5p�PJ��
�`V��a�z�58`RѡCM���r�MpR^pE��dQ_P�R�`�uMq���c$p�YSL�p�`� � q�'⏇��f����`0��"d��VALU���J����Q[hFaIgD_L�eHI~j�I��$FILE_q��d��$�j�c�SA+�� h � �VE_BLC�Kˣ�bj��hD_CPU yr� yfК��o��d�pYO�k�R � � PWR�����aqLA��S�*�fswqptRUN_FLG�uet�qpt�� �u�qet�qpuHk�|tx�ppt��TBC2��_� � (�B�p�M���;�� ��.�TDC�p��!�π��/��TH.�J��TV��R�4�ESERV�E!�w�.�w�3t���$$CLAk� ���h���O��O� ���զ�����׹�IR�TUAL����AA�VM_WRK 2� � �0  �5ȯ��'��J� J�	m�^���O��!�o�������]�Н�ܟl���)�1���B�S��� 1Ɖ�? <�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f��x��A�C1�AXL�MTÀ���Z�  d��IN����PRE_EXE��1����QAT��R�����IOCNV_�NUM�� ȶ�P��US��V�@�IO�_$� 1�P $�痑�����?���P�������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v������LARMRECOV ������[�LMDG �k�v��LM_IF k����5� G�Y�k�y�#��������ҿ�, 
  �χ���2�D�V�h����ANGTOL � � 	 A�   �Ϲ˟�PP�LICATIONg ?�������ArcTo�ol �� 
V�9.00P/03���y�
8834�0���F07�$�1�612������7DC3�y���N�oney�FR=Ay� 6Tݚ�P_ACTIVJ������UTO�MOD
����P�_CHGAPON�L� �OUP�LED 1k��� Y�]�o����CUREQ 1k�W  T�������	�������Ф���_ARC �Wel��AW����AWTOPK7�HKY����� ���Q�c�u������� ��������)� M_q����� ��%I[ m������� �/!/{/E/W/i/�/ �/�/�/�/�/�/�/? ?w?A?S?e?�?�?�? �?�?�?�?�?OOsO =OOOaOO�O�O�O�O �O�O�O__o_9_K_ ]_{_�_�_�_�_�_�_ �_�_oko5oGoYowo }o�o�o�o�o�o�o�o g1CUsy� ������	�c� -�?�Q�o�u�������0��Ϗ	��TO�������DO_CLEA�N)���`�NM  ��������П������_DSPDR3YRg�:�HI���@��b�t��������� ί����(�:���MAX��G� ��8�X�XG��T����PLUGGG�H�T�X�WPRC�B����Q�C���O��"���SEGF �B� �� �����b�tφϘϪ���LAP?�R�� ����(�:�L�^�p���ߔߦ߸��߿�TO�TALz���USE+NU?�L� -�1����RGDISPWMMCB�J�C�O�@@��L�O=��_�-�RG_STRING 1�
�M�S���
��_ITE;M1��  n���� ����	��-�?�Q�c� u����������������)I/O SIGNAL���Tryout� mode��I�npi Simul�ated��Ou�t{OVER�R<� = 100���In cyc�lo��Prog� Abor���~estatus��� cess Fa�ult�Aler��	Heartb�ea�KHand? Broke>; =Oas�����C���C���� ///A/S/e/w/�/�/ �/�/�/�/�/??+?p=?O?a?�WOR� ��1/s?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O_^PO��=P�;&_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono��o�o�o�o8RDEV @^�`T_�o,> Pbt����� ����(�:�L�^�PALT����? _�����я����� +�=�O�a�s�������ໟ͟ߟ�s�GRI ]���)����Q�c�u� ��������ϯ��� �)�;�M�_�q�������R�ͱA����� ��+�=�O�a�sυ� �ϩϻ���������x'�9߻�PREG�� r��Kߙ߽߫����� ����)�;�M�_�q��������?��$ARG_�0D �?	��� ���  w	$?	[4��]4��?U��SB�N_CONFIG� �srm�C�II_SAVE � ?����T�CELLSETU�P 
 �%  ?OME_IO??%MOV_H������REPм:�UTOBACK��� ���FRA;:\_� A_֖��'`� _׊� ��� �23/04/0�8 11:47:14_�V�_��	6-{��V}� ����_քk/ /)/;/M/_/��/�/ �/�/�/�/�/z/?%? 7?I?[?m?�/�?�?�?��?�?�?�?۰�  �v_Y_\ATB�CKCTL.TM�P DATE.D���DOVOhOzO�OSIKNI�����S?MESSAG��A���(�KODE_D ��������EO�`�O�SPAUS=Q!�� � ,,		��  �M_[WA_ {_e_�_�_�_�_�_�_ �_�_/ooSo=oOo�o��� T*PTSK � 0]��OV UP3DT�@�Gd�`�F�XWZD_ENB8�D��vSTA�E ���e�WEPLSC�H Rb   �fj|�� �������0� B�T�f�x��������� ҏ�����,�>�P�nDsROD,r2 ���Lڳ�� %��ɟ۟����#� 5�G�Y�k�}�������WEROBGRPƮh[r�b��WEWELn�������� ?�Q�c�u����������Ͽ����
�XI-Ss�UN� ���ա� 	�of�:�U� ��yϲϝ����������
�0�3�METERs 2�f�� P��t�ߘ�+�SCRD�CFG 1 ��l ����� ������'�9�K���Q���ߛ����� ����\����=�O�a��s�������8�KYG�R;��`_��@NA�ME 	�	�Y��_ED�@1���� 
 �%=-%@EDT-��#�Tx��� *�? G|�0��'�?������2�"�6 �GÕ}��l��3�%/I[��I/��8/��4 �/��//[�/?\/n/?�/�5M?�/�? �/[v?�?(?:?�?^?�6O�?fO�?[BO@�O�?O�O*O�7�O UO2_yO[_y_�O�Oh_�O�8�_Y�_}�\�_Eo�_�_4o�_B�9}o�_�oo�\��oXojo �o�CR� _��V]p��"4�X��# NO�_DEL����GE?_UNUSE�����IGALLOW �1�   (�*SYSTE�M*�	$SER�V_á|ٕ�POS7REG��$��|܎��NUMÊ�֍�PMUA��LA�YM�|�PM�PALT�CYC10"�5��#�[�ULSU�׍7�����Lq���BOX�ORIǅCUR_���֍PMCNV6���10K���?T4DLIB�����	*PROGRA���PG_MI#�M�_�AL-�l�V��_�B����$F�LUI_RESUP;�ï͏�s�|� �"�4�F�X�j�|��� ����Ŀֿ����� 0�B�T�f�xϊϜϮ� ����������,�>��P߳x��LAL_OUT �����WD_ABOR<��e���ITR_RT/N  �d�����?NONSTO ��� M�CCG_C�ONFIG  
����:ㆃD�R��E_RIA_Ib����z����F?CFG 
.�z�m��_LIM���2- <��# 	�����b<���j-���`���PA���GP 1�����i�{���L��C������C1��9���@���C��CV���]��d��l��s���d�C[��m���v���������� C���D �6�g?��HE�����]G_Pݐ15� -�P������\�HKoPAUS��1��z� K�(n��\ ������/� *//:/`/F/�/�/|/4�/X�O�����g���COLLECT�_����М�7E�N-�����2�!ND-E3��P��r�1234567890o7�b����m?�6�c
 Hy��c) �?�?�|�?�?$O�{�? OhO3OEOWO�O{O�O �O�O�O�O�O@___ /_�_S_e_w_�_�_�_ �_o�_�_o`o+oI6:��; ��I6IO !X91�h����o�o�gTR�0�2"�m(�`�i
Ao&~"�#�mPzn^�i_MOR��$5� �R	�u���y�����9�'��r+��%J�},n?WW���R�`K���aZR���&�/ŏāĂC4 W A����`x�`�A��Cz  B��C�0BO 	�C�  @���`^�a:d�
��IQ3�'����T_DE-Fx� l�%^y�<�M�INUS:�m�z厔KEY_TB�L  4�z�Ā� �	
��� !"#$%&'�()*+,-./�x7:;<=>?@�ABCP�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������S���͓���������������������������������耇���������������������9��a��LCK��露���STA�ߌ�_AUTO_DO�9���IND04 ��1R_T1��T�2Z�� �A���XC�*� 2(���08�
SONY XCg-56ɏÁࣀ_�@���1� Kp�А̵HR�5�9Ns���R57<�"�Aff.�h��ϖ� rϻ��Ϩ��� ���'�9��]�o�J���ߥ߀�����i|TR�LO�LETEo��J�T_SCREE�N 5�k�csc\U��MM�ENU 1)5�  <��g�� �^���#������ ����/���e�<�N� t������������� ��(a8J�n ������� K"4�Xj�� �����5/// D/}/T/f/�/�/�/�/ �/�/�/1???g?>? P?�?t?�?�?�?�?�? O�?OQO(O:O`O�O pO�O�O�O�O_�O�O�_M_$_6_�_ylA�_?MANUAL��Q��DBwq~r��DB�G_ERRLU�9*M��a �_o�*o<n�QNUML+IM��`d��,��DBPXWORK 1+M�o�o�o�o�o�og}DBTB_�� ,�]؃Hq�Ä�QDB_A�WAY�S�GC;P ��=��lb:r�_ALX` �6r�RYЕ�	开�X_�P 1�-��q|�
��o�Ȅ���h_M&7�IS��E{@����ONTIM��&���,��y
���sMOTNEND����tRECORD ;13M� ���sG�O����{Er � ��$���,�S� w�換�����V�l��� d����=�O�a�s�� �����*�߯��� ��9���]�̯������ ��&�ۿJ���n�#�5� G�Y�ȿ}�쿈���� ������j�ߎ�߲� g�yߋߝ���߬ߺ���f�f�-�?��c� N��ߙ��p�U���� ��[���4����wt� g�y���������B��|DJ_��-�� Q<J������>�TOLERE�NCCtBȌrQpL����PCSS_C�NSTCY 24Jzi��P��r�D Rdv����� ��//*/</N/d/�r/�/�/DEVI�CE 25/ v�/�/??1?C?�U?g?y?�?�?� HNDGD 6/�#pCz�>LS 27�-�?O-O?OQO�cOuO�O�?!PARAM 8�ysr�U��DSLAVE� 9�=�7_CF�G :�O�Cd�MC:\!L%04d.CSV�Ob�pc8_�RyA eSCHmP�1��Nx_�_�G��F�R�Q�_x�Y�QPJP��S�^�qq�LRC_?OUT ;�-q��O_SGN <�����Q08-�APR-23 11:48hPyo�c�& V�^�i��a�N�`��mE�@�S�Þ��j��a�n�CVERSION lj�V4.0.1� �EFLOGIC� 1=/ 	��XPPy�Q`}2rPROG_ENBw�\�6�sULS7� �6�2r_ACCLI�M8���C�~�sWRSTJN�0�偃Q2qMO�|�Q��B �INIT �>/��Q �vO;PT�@ ?	=���
 	R57Y5�Cj�74o�6p��7p�50��%t��2�p��X��,wM�TO C Y��o�-vV$��DEX�wd�r`�+�PATH AljA\�x�����HCP_CLNT�ID ?v�C �k�ʟ�IA�G_GRP 2C�
Y �� �	 D�  D��� D  Bu��ff�� �?���<��h��V���B�N��C�-Bz���Bpe`���mp2m7 7�89012345�6�����  �Ao�mAj�1AdA]��
AW|�AP���AJ-AC/A;�A4-�Lؠa@�eT��A��A�hPB�4��� ��Y�a
�עuƨApff�Aj�yAeK��A_�AY���ASy�MC�AF?��A@ �9���"�4�9�H�9�W�@��X�ȑ�@��y������ſ׿�鸃;d5?�@~ff@x1'�@q��@kC��@d�D@]��@Vv��-�?�Q��c��s��l��@�e@^��@�W\)@O��@�pP@?!�7K�@.V�Ϲ������Ͼ�S@M�G�!�A��@<1�@5��@/l��@(Ĝ@!���\3�E�W�i�{�]� �/�A��e�w��K� ������������ =�O�-�s������A� ��x�����Ѩ�/��>��R��?�3�3?Y����̽�/�7'Ŭ6� 4�F#���L/�@�p�?��
=@�@��Q�O�m@,�Ah�eP�eP�9�= c�<��]>*��H>V>�3��>���/�<���<� ���^� �?� �C�  <(�U�Rw 4;�33�X���	��A@�R?7� ��)��7]o;�� {�?����/޻�?�73!>��(�>��?!=�ʽ�/���G�[/G��/����Ռ%����|eP� @���@hP?@Q�?L�����ŗ�Iߟ5�˦(�G?�"��'�p%1�0?{&��L4V?5�C�>qP���C'^?�,��?�? <�P �?�?�?�T�?O�?=O�+[HgH��O &O�O�O�O�O�O_�O�%_�CT_CON�FIG D��|��deg�U��STBF_TTS�w
�ywSp�s�Q:�V/`MAU�p�~�rMSW_CFKP�E��  0�VjOCoVIEW�PF�]:���ޟ0oBoTofo xo�o�o�o�o�o�o �o�o1CUgy ������	� ��?�Q�c�u����� (���Ϗ������ ;�M�_�q�������6� ˟ݟ���%���I��[�m�������\RC�SGg��R!?���ۯ ���4�#�X�G�|��T�SBL_FAUL�T HΪ�X��G�PMSK�W��?PTDIAG IOY��Q�)UD1�: 678901�2345�\X=P _B�T�f�xϊϜϮ� ����������,�>�P�b��8 t:�
1Ϫ�9VTREC	P߿�
����?*� '�9�K�]�o���� �����������#�5��G��߀ߒߏ�2]UM�P_OPTION�P����TR�R�S�����PMEU��Y�_TEMP  ?È�3B��P$ s�A! UNI�P��U$ѶYN_BR�K J	o<RED�IT_��ENT �1KΩ  ,�&CL_DES�CARGAEPVEcYO�P�`&� �CAPTURA_?INDEX ���'&��X����FP��	IR_?A_HOME��?PLACE�w��9&PICK_Nw RAD�.�
�����l� /\R� �+//O/6/^/�/l/ �/�/�/�/�/?�/'? 9? ?]?D?�?h?z?�?�?�?�=m MGDI_STA7�Q$h�NCC1L�[ ��[�MO@O��
��d ���O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o�� 8oJo\ono|i�A|o�o �o�o�o�o�o 2 DVhz���� ���
��j1o;�M� _�q��o������ˏݏ ���%�7�I�[�m� �������ǟٟ��� �)�3�E�W�i����� ����ïկ����� /�A�S�e�w������� ��ѿ����!��=� O�a�{�qϗϩϻ��� ������'�9�K�]� o߁ߓߥ߷������� ���+�5�G�Y��� ������������� �1�C�U�g�y����� �����������#�- ?Qc}���� ���);M _q������ �/%/7/I/[/u /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?/O /OAOSOm/_O�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_O�_'o9oKoeO wO�o�o�o�o�o�o�o �o#5GYk} ������oo �1�C�U�ooy����� ����ӏ���	��-� ?�Q�c�u��������� ϟ�[���)�;�M� g�q���������˯ݯ ���%�7�I�[�m� �������ǿٿ�� �!�3�E�_�i�{ύ� �ϱ����������� /�A�S�e�w߉ߛ߭� �����������+�=� W�M�s������� ������'�9�K�]� o��������������� �#5��a�k} ������� 1CUgy�� �������	//-/ ?/Yc/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? �OO%O7OQ/[OmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�?�_oo /oIO;oeowo�o�o�o �o�o�o�o+= Oas����� �_���'�AoSo]� o���������ɏۏ� ���#�5�G�Y�k�}� ������ş����� �1�K�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� 7�����)�C�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ�������� �!�;�E�W�i�{�� ������������� /�A�S�e�w������� ��������3�) Oas����� ��'9K] o��������� �/�=G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?���?�?	OO5/ ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�?�_ �_oo-O7oIo[omo o�o�o�o�o�o�o�o !3EWi{� ���_����%o �A�S�e�w������� ��я�����+�=� O�a�s���������� ߟ���/�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������͟׿���� '�1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ��ſ ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� �!3EWi{� ������ /ASew���� ����/+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]?�o?�?�?� �$E�NETMODE �1M%��  ����?�;�0RROR�_PROG %��:%�/O<I
ETA�BLE  �;�/{O�O�O�G
BSE�V_NUM �2?  ��1�@�
A_AUTO_ENB  �5�3Dw_NO�A N�;��1�B  *�*'P�'P�'P�'P�@�+&P@_R_d_ THI�S�C��0�K_AL�M 1O�; �2�'\�+e_�_@�_oo)o;oi__�B.P  �;%Q�2��j�0TCP_VE/R !�:!'OKo�$EXTLOG_7REQ�V��I�c�SIZ�o�dSTK��iU��bTOoL  �Dz�R��A �d_BW�D``5p�Faq�2JsD�IOq P%�es�4�f{STE�Pw��0�pOP_�DO�1FACTORY_TUN�W�d�yDR_GRP� 1Q�9�Ad 	�{o9��0*��*u����RHB� ��2 ���� �e9 ��� m�*����z�����׏ ����
��U�@��y�d�@ec5A?�@F�s���
 B�|�� �����8zc�j�����3��B�  Q�Aݠ���33]��3�3�@UUTy�@𗐊���7>u.��>*��<������E�� F@� ɢ�5Wե��J���NJk�I�'PKHu��IP�sF!�����?�  ���9��<9�8�96C'6<�,5������L{��1"���ZT6p� m�ߵ�l�jBKFE�ATURE R�%ap�1ArcTool ����Engli�sh Dicti�onary��4D� Standar�d��Analog� I/O��Aɰe� Shift�r�c EQ Pro�gram Sel�ect1�Soft�par&�1�Wel�d>�cedureys/ɯ�Core`����Rampingn�utoW�wa���Update��m�atic Bac�kup����gro�und Edit�����Cameraz�F
�Cell���nrRndIm���&�ommon �calib UI�!�e�sh5�]ߋ�c��ĝ�Y�ne����t%y�sH�c�n�p�Monitor���ntr��eliayb���DHCP���&�ata Acq�uis��%�iag�nos���?�oc�ument Vigewe�'�ua���heck Saf�etyx���han�|� RobF�rvB�q��yս���s���FC�����xt w�eav��ch��x�t. DIO��nsfi���end��Err�Lt�A���%s@�r�0� Pp���FCTN Men�u�����TP I�n��fac����G�en�ls�Eq �Lv����p Ma�sk Exc��g��HT��?�xy �Sv��igh-wSpe��SkiX��m���mmuni�c��on��Hou�r����:����co�nn��2rncr���struҲ��K�AREL Cmd7. L��ua��Run-Ti�E�nv�����+��s���S/W��Lic�ense���W�B�ook(Syst�em)��MACR�Os,2/Off;se��MMR����s�MechStoEp>�tJ�Y�9iR�"ˍx������od �wit�����h�.���Optm8�a?�fil��`�gh9ulti-�T��ƿ�PCM 'fun�i)oV�⼴ĉ-Regi.r,��l&ri��Fy+�&��NuE�Y��(C�AdjuF �.C�#�=tatu�!-?�����RDM��otϰs�coveرi5em�4�n�i5u2��	N��uesLŨ7o������SNPX b����SN��Cli���>#���r׳O�Q ����5ot��ssag���5.����?�` ��QzN/I|���EMILIB�O~�BP Firm��:�NP��Acc�
��TPTX4�Del�nQ�O�A��M�Mo�r�0 SimulQa��EVu�P���|J�!��&>�ev�.�E��ri��_?USB po^�p��iPK�a���Unexcept���0�$X�U����VCt�rQH�VU�6b�OGeK�AkS�0SCUyoS�UI��W�b(�lb PlD6�n��h�d  ���w�t�|6 ux�V�oCwGridy1play=}�@��Ww�R-b.�9-10�iA/7LMA�larm Cau�se/�0edٸA�scii>�Loa9d���zUpl�p��l˰��Gu��/�P���yc��� �P����RA�PC��i���`��l�p3c���NRT�z��Online HelX��m&��l&� �!�qtr���64MB DRsAM���FRO(��Z�t� .��ma�i��KŅL�Su�p�R*!�)��K���c�roE<t3E�tAfrt��t3���<����� �=�4�F�s�j�|��� ����̯֯����9� 0�B�o�f�x������� ȿҿ�����5�,�>� k�b�tϡϘϪ����� �����1�(�:�g�^� pߝߔߦ���������  �-�$�6�c�Z�l�� ������������)�  �2�_�V�h������� ����������%. [Rd����� ���!*WN `������� �//&/S/J/\/�/ �/�/�/�/�/�/�/? ?"?O?F?X?�?|?�? �?�?�?�?�?OOO KOBOTO�OxO�O�O�O �O�O�O___G_>_ P_}_t_�_�_�_�_�_ �_oooCo:oLoyo po�o�o�o�o�o�o	  ?6Hul~ �������� ;�2�D�q�h�z����� ˏԏ���
�7�.� @�m�d�v�����ǟ�� П�����3�*�<�i� `�r�����ï��̯�� ��/�&�8�e�\�n� ��������ȿ����� +�"�4�a�X�jτώ� �ϲ���������'�� 0�]�T�f߀ߊ߷߮� ��������#��,�Y� P�b�|������� ������(�U�L�^� x��������������� $QHZt~ ������  MDVpz�� ����/
//I/ @/R/l/v/�/�/�/�/ �/�/???E?<?N? h?r?�?�?�?�?�?�? OOOAO8OJOdOnO �O�O�O�O�O�O_�O _=_4_F_`_j_�_�_ �_�_�_�_o�_o9o 0oBo\ofo�o�o�o�o �o�o�o�o5,> Xb������ ���1�(�:�T�^� ����������ʏ���  �-�$�6�P�Z���~� ������Ɵ����)�  �2�L�V���z����� ��¯����%��.� H�R��v��������� ����!��*�D�N� {�rτϱϨϺ����� ����&�@�J�w�n� �߭ߤ߶�������� �"�<�F�s�j�|�� ������������ 8�B�o�f�x������� ������4> kbt����� �0:g^ p������	/  //,/6/c/Z/l/�/ �/�/�/�/�/?�/?�(?2?_?V?h?�?  �  H5�41�3�12�6R7�82�750�5J6�14�776�5AW�SP�71�7RCR��88�6TU�6J5�45�8�6VCAM޴5CLIOPFRI�OGUIF�666GC�MSC�H�6STY�L�72FCNREv�652�6R63�7�SCH�5DOCV��FCSU�5ORS^FR869�70�7�88�6EIO�FR�54�6R69�6E�SET,GGJIW{MG�5MASK�5�PRXY�H7�6O	C[F`P3,H�6`P�8��853VH�XLC�H�VOPL{VJ5m0�VPS
gMC�7�`cW55�6MDS�WHg�WOP�WMP�R[F�@�VP�6PC�MsG0�g`P�750��g517G51�h0n7FPRSWW69�V�FRDOFRMCNܘFXH93�6SN�BAtG�WSHLBb�FMNw�@�GNN�X�2�6HTC�6TMqI�F�0VTPA�FoTPTX�vELv�`W8�7�0�6J9�5FTUT�W95�VUEC�VUFR�OFVCC'�OFV;IP�FCSC�v�@�Ih�6WEB�6H�TT�76�GWIO�c�CG��IGb�I�PGS��RC�FH�77�7667FR7�JWR�hR53�88j�h2�VR�Y64W54��66�6|@�6�NVDWVD0R�Fnu�CTO+GNN�V�OL�HEND�6L2�FVR�E�8ҟ� ����,�>�P�b�t� ��������ί��� �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D� V�h�zߌߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N�`�r��� ������������ &8J\n��� �����"4 FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/??,?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O �O�O�O�O�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�o�o�o �o�o
.@Rd v������� ��*�<�N�`�r��� ������̏ޏ���� &�8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�������į ֯�����0�B�T��f�x�����  ?H541�����2��R782��5�0��J614�7�6��AWSPȻ1��RCR��8�T=U�J545���VCAM��CLI�O��RI��UIFzȺ6f�CMSC��^�STYL�2G�oCNREȺ52�wR63ǻSCH���DOCVH�CSUORS7�R86�9�0��88��E�IO��R54׺R{69�ESETX˺&�J%�WMG��M�ASK��PRXY���7��OC����3`X�׺����53���H��LCH'�OP�L�J50g�PS���MC�����55���MDSW(�V�OPV�MPR��4�G�\���PCM��0��l����50w�51g��51��0g�PRSv��69G�FRD���RMCN��u�H9=3�SNBA�ˆ�/SHLB��M�4��'�NN��2�HTC�TMI��԰���TPA��TPTXF�
EL7
����8ֻ�԰��J95G�TU�TW�95G�UEC�'�UFR��VCC��O7�VIP��C�SCe�I����W�EB�HTT�6n&�WIO�CG&+{IG�IPGSX*�RC��H77ǻ6�6g�R7��R��R�53��8��2g�R���64��54�+6q6������NVD���D06;Fe<CTO�W�NNG�OL��E�NDȺL�FVR �ɗ��?�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H��Z�l�~������STD��LANG����Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas�p����RBT��OPTN��p,>PbDPN�� z�������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ ޟ���&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ���� �0�B�T�f�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\?�n?�?�:99�5��$FEAT_AD�D ?	�����1�0  	�8�?�?�?
OO.O @OROdOvO�O�O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|� �������� 0�B�T�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�\�n�����������4DEM�O R�9   �8����2 );h_q��� ����.%7 d[m����� ���*/!/3/`/W/ i/�/�/�/�/�/�/�/ �/&??/?\?S?e?�? �?�?�?�?�?�?�?"O O+OXOOOaO�O�O�O �O�O�O�O�O__'_ T_K_]_�_�_�_�_�_ �_�_�_oo#oPoGo Yo�o}o�o�o�o�o�o �oLCU� y������� 	��H�?�Q�~�u��� ����؏Ϗ���� D�;�M�z�q������� ԟ˟ݟ
���@�7� I�v�m������Яǯ ٯ����<�3�E�r� i�{�����̿ÿտ� ���8�/�A�n�e�w� �ϛ��Ͽ�������� 4�+�=�j�a�sߍߗ� �߻��������0�'� 9�f�]�o������ ��������,�#�5�b� Y�k������������� ����(1^Ug �������� $-ZQc}� ������ // )/V/M/_/y/�/�/�/ �/�/�/�/??%?R? I?[?u??�?�?�?�? �?�?OO!ONOEOWO qO{O�O�O�O�O�O�O ___J_A_S_m_w_ �_�_�_�_�_�_oo oFo=oOoioso�o�o �o�o�o�oB 9Keo���� �����>�5�G� a�k�������Ώŏ׏ ����:�1�C�]�g� ������ʟ��ӟ ��� 	�6�-�?�Y�c����� ��Ư��ϯ����2� )�;�U�_�������¿ ��˿����.�%�7� Q�[ψ�ϑϾϵ��� ������*�!�3�M�W� ��{ߍߺ߱������� ��&��/�I�S��w� �����������"� �+�E�O�|�s����� ����������' AKxo���� ���#=G tk}����� �///9/C/p/g/ y/�/�/�/�/�/�/? 	??5???l?c?u?�? �?�?�?�?�?OOO 1O;OhO_OqO�O�O�O �O�O�O
___-_7_ d_[_m_�_�_�_�_�_ �_o�_o)o3o`oWo io�o�o�o�o�o�o �o%/\Se� �������� !�+�X�O�a������� ď��͏�����'� T�K�]����������� ɟ������#�P�G� Y���}�������ů� �����L�C�U��� y������������� ��H�?�Q�~�uχ� �ϫϽ��������� D�;�M�z�q߃߰ߧ� ��������	��@�7� I�v�m������� ������<�3�E�r� i�{������������� 8/Anew ������� 4+=jas�� �����/0/'/ 9/f/]/o/�/�/�/�/ �/�/�/�/,?#?5?b? Y?k?�?�?�?�?�?�? �?�?(OO1O^OUOgO �O�O�O�O�O�O�O�O $__-_Z_Q_c_�_�_ �_�_�_�_�_�_ oo )oVoMo_o�o�o�o�o �o�o�o�o%R I[�����}  �x�	� �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q��������� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s��������������   ������1CU gy������ �	-?Qcu �������/ /)/;/M/_/q/�/�/ �/�/�/�/�/??%? 7?I?[?m??�?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{�����������
��������# 5GYk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{�������y�$FEAT�_DEMOIN [ �t����p}�tINDEX�����pILEC�OMP S�;��M���u�C�SETUP2 �TM�W���  N ��@�_A�P2BCK 1U~M�  �)�xD��ŋ%����pP� ׏��u��@�Ϗd�� q���)���M������ ���<�N�ݟr���� ��7�̯[�����&� ��J�ٯn������3� ȿڿi�����"�4�ÿ X��|�ωϲ�A��� e���ߛ�0߿�T�f� �ϊ�߮���O���s� ���>���b��߆� ��'��K������� ��:�L���p����#� ����Y���}�$�� H��l~�1� �g�� �-V �z	��?�c �
/�./�R/d/� �//�/;/�/�/\����P�� 2��*�.VR�/3?� *�6?\?�#b?�?p%0P�C�?�?� FR6�:�?�>r?O�;T +�+O=O�5(OgL��?<�Oo&*.F ?�O"�!	�3�O�LzO_�KSTM_D_�2�0D0_o]�O�_�KH`_��_UW�_q_�_o�JGIF"oLoWU8o�_o�o�JJPG�o�oWU`�oyo�o �:JS*�S� �cA�o%
�JavaScri3pt�oCSp��VV�� %Ca�scading �Style Sh�eets�u 
A�RGNAME.D)T2��,ZP\F���fqv���3�v�DISP*}�`�ZPʏ
�������
TPEINS.XML:���:\N��n�Cu�stom Too�lbar����PA?SSWORD��.?FRS:\ҟ��� %Passw�ord Config�n/\��U��� �/��E�گ�{���� 4�F�կj������/� ĿS��w��ϭ�B� ѿf�x�Ϝ�+����� a��υ�ߩϻ�P��� t��mߪ�9���]��� ��(��L�^��߂� ��5�G���k� ��� ��6���Z���~���� ��C�����y���2 ����h����� Q�u
�@� dv�)�M_ ��/�/N/�r/ /�/�/7/�/[/�/? �/&?�/J?�/�/�?? �?3?�?�?i?�?�?"O 4O�?XO�?|O�OO�O AO�OeOwO_�O0_�O )_f_�O�__�_�_O_ �_s_oo�_>o�_bo �_o�o'o�oKo�o�o �o�o:L�op�o ��5�Y�}� $��H��A�~���� 1�Ə؏g����� �2� ��V��z�	����?� ԟc�͟
���.���R� d�󟈯�����M�� q������<�˯`�� Y���%���I�޿�� ϣ�8�J�ٿn������!�3��ϫ��$FI�LE_DGBCK� 1U������� <� �)
SUMM?ARY.DG��~�OMD:�F����Diag Su�mmaryG�T�
CONSLOG<���1ъ���Y�Co�nsole lo�g��S�	TPACCN��%�%�J�U��TP Acco�untin��T��FR6:IPKD?MP.ZIP~���
����V�f�Exc?eption����2�MEMCHEC�K@��5�V���M�emory Da�taW���+YF)	FTP�߮�=����a���mmen�t TBD����L� =�)ETHERNET��|���^Y�Ethe�rnet ��fi�gura��Z���DCSVRF��������g�%�  v�erify alyl���M+��DIFF���e�h�%�dif�fg� CHG01\CU��},/*f�2��@�n/y/!/�3d/8K/]/�/ �/?��&VTRNDIAG.LS?�/�/�v?i�61 ^�no�sticw?��T6�a)UPDA�TES.�0�?��FRS:\�?�=�Z�Updates� List�?|�P�SRBWLD.C	M*O~��2>O�?���PS_ROBOW�EL��R�b1HADOWl?Q?c? _g��Shadow Changes_��q�BNOT�I��O�O�_e�N?otific�'_��+@AG`��_�� �_��
o3oZ�Wo�_{o �oo�o@o�o�ovo �o/A�oe�o� ��N�r��� =��a�s����&��� ͏\�񏀏���"�K� ڏo�������4�ɟX� �����#���G�Y�� }����0���ׯf��� ���1���U��y��� ���>�ӿ�t�	Ϙ� -ϼ�:�c���ϫ� ��L���p��ߦ�;� ��_�q� ߕ�$߹�H� ����~���7�I��� m��ߑ��2���V��� ���!���E���R�{� 
���.�����d����� /��S��w� �<�`��+ �Oa���� J�n//�9/� ]/�j/�/"/�/F/�/ �/|/?�/5?G?�/k? �/�?�?0?�?T?�?x? �?O�?CO�?gOyOO �O,O�O�ObO�O�O_ -_�OQ_�Ou__�_�_ :_�_^_�_o�_)o�_ Mo_o�_�oo�o�oHo �olo�o7�o[ �o� �D�� z��3�E��i�� �����ÏR��v�� ���A�Џe�w���� *���џ`�������� &�O�ޟs������8� ͯ\�����'���K� ]�쯁����4���ۿ����$FILE_�FRSPRT  ���Ű�����MDO?NLY 1UŽ�� 
 �)�MD:_VDAEXTP.ZZZ����j�y�6%�NO Back �file DϽ�S�6p���Z��ϸ� ��%�j�I���m��� ��2�����h��ߌ�!� 3���W���{�
��� @���d������/��� S�e���������N� ��r���=��a ����&�J�����9K��VI�SBCK"��1��*.VDL��FR:\eION?\DATA\�'�Vision VD����
/ /2@/*d/�u/�/ )/�/M/�/�/�/?�/ <?�/�/r??�?�?c? �?[?�??O&O�?JO �?nO�OO�O3O�OWO iO�O�O"_4_�OX_�O |__�_�_A_�_e_�_ o�_0o�_To�_�_�o��LUI_CON�FIG V��x�k $ sc'�{��o�o"04FTy�`|x|o~ �����|l�� �/�A��R�w����� ����V������+� =�ԏa�s��������� R�ߟ���'�9�П ]�o���������N�ۯ ����#�5�̯Y�k� }�������J�׿��� ��1�ȿU�g�yϋ� ��4Ϯ�������	�� ��?�Q�c�u߇ߙ�0� �����������;� M�_�q���,���� ��������7�I�[� m����(��������� ����3EWi{ �$������ 
/ASew� ������/+/ =/O/a/s/
/�/�/�/ �/�/�/�/?'?9?K? ]?o??�?�?�?�?�? �?�?O#O5OGOYOkO O�O�O�O�O�O�O�O __1_C_U_�Of_�_ �_�_�_�_j_�_	oo -o?oQo�_uo�o�o�o �o�ofo�o); M�oq����� b���%�7�I�� m��������ǏZ��@���!�3�E�Ոa��|�$FLUI_�DATA W����v��فh�RESUL�T 2Xv���� �T�/w�izard/gu�ided/ste�ps/ExpertQ�֟�����0��B�T�f�x�������Continue with G��ance��ӯ��� 	��-�?�Q�c�u����� _�-`�v���0 �း�x�lw�ع���ps�� #�5�G�Y�k�}Ϗϡ� �������Ϩ���"� 4�F�X�j�|ߎߠ߲� ��������ؿʿܿ�}��torch� p�����������  ��$�6���Z�l�~� ��������������  2D��_9�K�wproc_��� ��0BTf x�I������ //,/>/P/b/t/�/@�/Wi�/��������TimeUS/DST�/*?<?N?`? r?�?�?�?�?�?�?��Disabl�� O%O7OIO[OmOO�O��O�O�O�O�N_�ـ�/�/�/�/�/224?z_�_�_�_�_ �_�_�_
oo.o�?�? dovo�o�o�o�o�o�o �o*<�O__�1_󷩟��Region?������(�:�L�^�p�����America� ��Ώ�����(�:�@L�^�p�����Jqy���j̟��
2Edi Z���"�4�F�X�j�|��������į֯� T�ouch Pan�el � (re�commen	�) �)�;�M�_�q����� ����˿ݿ�������� ����
2acces��uχϙϫϽ����������)ߘC�onnect t�o Network8�o߁ߓߥ߷��߀�������#�5�0X�t�6��!J�0�Introduct���������'� 9�K�]�o�������� ��������#5G0Yk}� �/b� ���HR��&8 J\n����� ����/"/4/F/X/ j/|/�/�/�/�/�/Fx�� ��
���~ ?*?�Q?c?u?�? �?�?�?�?�?�?OO )O�MO_OqO�O�O�O �O�O�O�O__%_�/ �/??|_>?�_�_�_ �_�_�_o!o3oEoWo io{o:O�o�o�o�o�o �o/ASew �H_Z_l_��_�� �+�=�O�a�s����� ����͏�o���'� 9�K�]�o��������� ɟ۟��� ��G� Y�k�}�������ůׯ �����ޏ0�U�g� y���������ӿ��� 	��-��N��r�4� �ϫϽ��������� )�;�M�_�q߃ߔϧ� ����������%�7� I�[�m��>Ϡ�b��� �������!�3�E�W� i�{������������� ��/ASew ���������� ���Oas�� �����//'/ ��K/]/o/�/�/�/�/ �/�/�/�/?#?�D? h?z?>/�?�?�?�? �?�?OO1OCOUOgO yO8/�O�O�O�O�O�O 	__-_?_Q_c_u_4? ~?X?�_�_�?�_oo )o;oMo_oqo�o�o�o �o�o�O�o%7 I[m���� �_�_�_���_E�W� i�{�������ÏՏ� �����oA�S�e�w� ��������џ���� �����p�2��� ����ͯ߯���'� 9�K�]�o�.������� ɿۿ����#�5�G� Y�k�}�<�N�`��τ� ������1�C�U�g� yߋߝ߯��߀����� 	��-�?�Q�c�u�� ������Ϡϲ�� ��;�M�_�q������� ����������$ I[m���� ���!��B� f(������� �////A/S/e/w/ ��/�/�/�/�/�/? ?+?=?O?a?s?2�? V�?z�?�?OO'O 9OKO]OoO�O�O�O�O �O�/�O�O_#_5_G_ Y_k_}_�_�_�_�_�? �_�?
o�?�_CoUogo yo�o�o�o�o�o�o�o 	�O?Qcu� �������� �_8��_\�n�2���� ��ˏݏ���%�7� I�[�m�,������ǟ ٟ����!�3�E�W� i�(�r�L�������� ����/�A�S�e�w� ��������~����� �+�=�O�a�sυϗ� �ϻ�z�į�����ԯ 9�K�]�o߁ߓߥ߷� ���������п5�G� Y�k�}�������� ������������d� &ߋ������������� 	-?Qc"� ������ );M_q0�B�T� �x���//%/7/ I/[/m//�/�/�/t �/�/�/?!?3?E?W? i?{?�?�?�?�?�� �O�/OAOSOeOwO �O�O�O�O�O�O�O_ �/_=_O_a_s_�_�_ �_�_�_�_�_oo�? 6o�?ZoO�o�o�o�o �o�o�o�o#5G Yk|o����� ����1�C�U�g� &o��Jo��noӏ��� 	��-�?�Q�c�u��� ������|���� )�;�M�_�q������� ��x�گ������¯7� I�[�m��������ǿ ٿ����Ο3�E�W� i�{ύϟϱ������� ���ʯ,��P�b�&� �ߛ߭߿�������� �+�=�O�a� υ�� �����������'� 9�K�]��f�@ߊ��� v�������#5G Yk}���r�� ��1CUg y���n������ /��-/?/Q/c/u/�/ �/�/�/�/�/�/?� )?;?M?_?q?�?�?�? �?�?�?�?O��� �XO/O�O�O�O�O �O�O�O_!_3_E_W_ ?{_�_�_�_�_�_�_ �_oo/oAoSoeo$O 6OHO�olO�o�o�o +=Oas�� �h_�����'� 9�K�]�o��������� vo�o�o���o#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	�ȏ*��N��u��� ������Ͽ���� )�;�M�_�p��ϕϧ� ����������%�7� I�[��|�>���b��� �������!�3�E�W� i�{����p����� ����/�A�S�e�w� ������l��������� ��+=Oas�� �������' 9K]o���� ������ /��D/ V/}/�/�/�/�/�/ �/�/??1?C?U? y?�?�?�?�?�?�?�? 	OO-O?OQO/Z/4/ ~O�Oj/�O�O�O__ )_;_M___q_�_�_�_ f?�_�_�_oo%o7o Io[omoo�o�obO�O �O�o�o�O!3EW i{������ ��_�/�A�S�e�w� ��������я����o �o�o�oL�s����� ����͟ߟ���'� 9�K�
�o��������� ɯۯ����#�5�G� Y��*�<���`�ſ׿ �����1�C�U�g� yϋϝ�\��������� 	��-�?�Q�c�u߇� �߫�j�|����߲�� )�;�M�_�q���� ��������� �%�7� I�[�m���������� ����������B� i{������ �/ASdw �������/ /+/=/O/p/2�/ V�/�/�/�/??'? 9?K?]?o?�?�?�?d �?�?�?�?O#O5OGO YOkO}O�O�O`/�O�/ �O�/�O_1_C_U_g_ y_�_�_�_�_�_�_�_ �?o-o?oQocouo�o �o�o�o�o�o�o�O �O8Joq��� ������%�7� I�om��������Ǐ ُ����!�3�E� N(r���^ß՟� ����/�A�S�e�w� ����Z���ѯ���� �+�=�O�a�s����� V���z�Ŀ��'� 9�K�]�oρϓϥϷ� �����Ϭ��#�5�G� Y�k�}ߏߡ߳����� �ߨ���̿޿@��g� y������������ 	��-�?���c�u��� ������������ );M��0�T� ����%7 I[m�P��� ���/!/3/E/W/ i/{/�/�/^p��/ �??/?A?S?e?w? �?�?�?�?�?�?��? O+O=OOOaOsO�O�O �O�O�O�O�O�/_�/ 6_�/]_o_�_�_�_�_ �_�_�_�_o#o5oGo X_ko}o�o�o�o�o�o �o�o1C_d &_�J_����� 	��-�?�Q�c�u��� ��Xo��Ϗ���� )�;�M�_�q�����T ��xڟ����%�7� I�[�m��������ǯ ٯ믪��!�3�E�W� i�{�������ÿտ� ���ʟ,�>��e�w� �ϛϭϿ�������� �+�=���a�s߅ߗ� �߻���������'� 9���B��f��RϷ� ���������#�5�G� Y�k�}���N߳����� ����1CUg y�J��n���� 	-?Qcu� �������// )/;/M/_/q/�/�/�/ �/�/�/����4? �[?m??�?�?�?�? �?�?�?O!O3O�WO iO{O�O�O�O�O�O�O �O__/_A_ ??$? �_H?�_�_�_�_�_o o+o=oOoaoso�oDO �o�o�o�o�o' 9K]o��R_d_ v_��_��#�5�G� Y�k�}�������ŏ׏ �o���1�C�U�g� y���������ӟ埤 ��*��Q�c�u��� ������ϯ���� )�;�L�_�q������� ��˿ݿ���%�7� ��X��|�>��ϵ��� �������!�3�E�W� i�{ߍ�L��������� ����/�A�S�e�w� ��HϪ�l���ϒ�� �+�=�O�a�s����� ����������' 9K]o���� ������� 2�� Yk}����� ��//1/��U/g/ y/�/�/�/�/�/�/�/ 	??-?�6Z?�? F�?�?�?�?�?OO )O;OMO_OqO�OB/�O �O�O�O�O__%_7_ I_[_m__>?�?b?�_ �_�?�_o!o3oEoWo io{o�o�o�o�o�o�O �o/ASew ������_�_�_ �_(��_O�a�s����� ����͏ߏ���'� �oK�]�o��������� ɟ۟����#�5�� ��z�<�����ůׯ �����1�C�U�g� y�8�������ӿ��� 	��-�?�Q�c�uχ� F�X�j��ώ����� )�;�M�_�q߃ߕߧ� ���ߊ�����%�7� I�[�m������� ���������E�W� i�{������������� ��/@�Sew ������� +��L�p2�� �����//'/ 9/K/]/o/�/@�/�/ �/�/�/�/?#?5?G? Y?k?}?<�?`�?� �?�?OO1OCOUOgO yO�O�O�O�O�O�/�O 	__-_?_Q_c_u_�_ �_�_�_�_�?�_�?o &o�OMo_oqo�o�o�o �o�o�o�o%�O I[m���� ����!��_*oo N�x�:o����ÏՏ� ����/�A�S�e�w� 6������џ���� �+�=�O�a�s�2�|� V���ʯ�����'� 9�K�]�o��������� ɿ������#�5�G� Y�k�}Ϗϡϳ��τ� �������ޯC�U�g� yߋߝ߯��������� 	��ڿ?�Q�c�u�� ������������ )������n�0ߕ��� ��������%7 I[m,���� ���!3EW i{:�L�^����� �////A/S/e/w/ �/�/�/�/~�/�/? ?+?=?O?a?s?�?�? �?�?�?��?�O� 9OKO]OoO�O�O�O�O �O�O�O�O_#_4OG_ Y_k_}_�_�_�_�_�_ �_�_oo�?@oOdo &O�o�o�o�o�o�o�o 	-?Qcu4_ �������� )�;�M�_�q�0o��To ��xoz����%�7� I�[�m��������ǟ �����!�3�E�W� i�{�������ï��� ����ޟA�S�e�w� ��������ѿ���� �؟=�O�a�sυϗ� �ϻ���������ԯ ���B�l�.��ߥ߷� ���������#�5�G� Y�k�*Ϗ������� ������1�C�U�g� &�p�Jߔ��������� 	-?Qcu� ���|��� );M_q��� �x�������/��7/ I/[/m//�/�/�/�/ �/�/�/?�3?E?W? i?{?�?�?�?�?�?�? �?OO�� /bO$/ �O�O�O�O�O�O�O_ _+_=_O_a_ ?�_�_ �_�_�_�_�_oo'o 9oKo]ooo.O@ORO�o vO�o�o�o#5G Yk}���r_� ����1�C�U�g� y����������o⏤o ��o-�?�Q�c�u��� ������ϟ���� (�;�M�_�q������� ��˯ݯ���ҏ4� ��X���������ǿ ٿ����!�3�E�W� i�(��ϟϱ������� ����/�A�S�e�$� ��H���l�n������ �+�=�O�a�s��� ���z�������'� 9�K�]�o��������� v���������5G Yk}����� ����1CUg y������� 	/����6/`/"�/ �/�/�/�/�/�/?? )?;?M?_?�?�?�? �?�?�?�?OO%O7O IO[O/d/>/�O�Ot/ �O�O�O_!_3_E_W_ i_{_�_�_�_p?�_�_ �_oo/oAoSoeowo �o�o�olO~O�O�O �O+=Oas�� �������_'� 9�K�]�o��������� ɏۏ�����o�o�o V�}�������şן �����1�C�U�� y���������ӯ��� 	��-�?�Q�c�"�4� F���j�Ͽ���� )�;�M�_�qσϕϧ� f���������%�7� I�[�m�ߑߣߵ�t� �ߘ��߼�!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� ��(��L�s�� �����' 9K]����� ����/#/5/G/ Y/z/<�/`b/�/ �/�/??1?C?U?g? y?�?�?�?n�?�?�? 	OO-O?OQOcOuO�O �O�Oj/�O�/�O_�? )_;_M___q_�_�_�_ �_�_�_�_o�?%o7o Io[omoo�o�o�o�o �o�o�o�O_�O*T _{������ ���/�A�S�ow� ��������я���� �+�=�O�X2|� ��h͟ߟ���'� 9�K�]�o�������d� ɯۯ����#�5�G� Y�k�}�����`�r��� �������1�C�U�g� yϋϝϯ��������� ���-�?�Q�c�u߇� �߽߫��������Ŀ ֿ�J��q���� ����������%�7� I��m���������� ������!3EW �(�:�^���� �/ASew ��Z�����/ /+/=/O/a/s/�/�/ �/h�/��/�?'? 9?K?]?o?�?�?�?�? �?�?�?�??#O5OGO YOkO}O�O�O�O�O�O �O�O�/_�/@_?g_ y_�_�_�_�_�_�_�_ 	oo-o?oQoOuo�o �o�o�o�o�o�o );M_n0_�T_ V�����%�7� I�[�m������boǏ ُ����!�3�E�W� i�{�����^���� �����/�A�S�e�w� ��������ѯ����� �+�=�O�a�s����� ����Ϳ߿񿰟��ԟ �H�
�oρϓϥϷ� ���������#�5�G� �k�}ߏߡ߳����� ������1�C��L� &�p��\��������� 	��-�?�Q�c�u��� ��X߽������� );M_q��T� f�x�����%7 I[m���� ����/!/3/E/W/ i/{/�/�/�/�/�/�/ �/���>? e?w? �?�?�?�?�?�?�?O O+O=O�aOsO�O�O �O�O�O�O�O__'_ 9_K_
??.?�_R?�_ �_�_�_�_o#o5oGo Yoko}o�oNO�o�o�o �o�o1CUg y��\_��_��_ 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ��4� �[�m��������ǯ ٯ����!�3�E�� i�{�������ÿտ� ����/�A� �b�$� ��H�JϿ�������� �+�=�O�a�s߅ߗ� V�����������'� 9�K�]�o���Rϴ� v�������#�5�G� Y�k�}����������� ����1CUg y�������� ����<��cu� ������// )/;/��_/q/�/�/�/ �/�/�/�/??%?7?��@d?�?�1�$�FMR2_GRP� 1Y�5�� �C4 w B�N 	 N ��?�<�0E�� �F@ �2�5W�EF:�0J��NJ�k�I'PKH�u��IP�sF�!��M?�  �JOF<�09�<9��896�C'6<,5���MA�  l�O�KBH�3B��0��@�A@�33�B�33F<�4�O]�0/@UUTZ@�@+P�MJ)>u.�>*���<���M=�[�B=���=�|	<�K�<�q�=�mbN���8�x	7�H<8�^6�Hc7��x2_ �__�_�_�_o o9o�L'�2_CFG =Z�;T Do�o��o�oKkNO ^�:
F0�a �`�JlRM_CHKTYP  �1N �0��0u0�1ROM�`_�MIN pN#���,p��@X�0SSB�[c[�5 �6YN%Psy��QeTP_DEF_�O@N$�3�wI�RCOM�`��$�GENOVRD_�DO!vW!�}TH�R!v d�ud�t_�ENB� �pRWAVC�3\BwMp� ��5Fs  �G!� GɃ��I�C�I(i J���ou���s�0"pÅF�G� �D�OU�0b��<�a�8���4<)p ^M6����.�P�~�N#C��0��0Ȕ�Sӟ��Ŗ���ē�9!��E�SM�T�3cR��0Op����$HOSTC[b1�d�9Np�W/ 5	y�y�y�L&��J)eů��� �,�:��]�o����������J�	anonymoul�ؿ��� � �2�x�����yϰ� үL���������>�� -�?�Q�c߆ϼ�ο�� ��������:�L�^�p� r�_�σ������ �����%�7�Z�� ������������ � 2�F�3z�Wi{ ������� d�ASew��� �����</+/ =/O/a/��/�/�/�/ �/�&8?'?9?K? ]?���v?�/�?/ �?�?O#O5O�?YOkO }O�O�?�O�/�O�O�O __f?x?�?�?y_�O �?�_�_�_�_�_>Oo -o?oQoco�_�O�O�o �o�o�o�o:_L_^_p_ ro_�_����� o���%�H6��o�m��������"�[�E�NT 1e� sP!I��  *���2�!�V��z�=� ��a�����ӟ����� ߟ@��d�'���K�]� ����⯥��ɯ*�� ��`�#���G���k�̿ ��ſ��&��J�� n�1�z�Uϣ��ϋ��� �����4���X��-����Q߲�u��ߙ�QUICC0�߿���2���13��!�����2��_�q���!ROUTER������"�!PCJOG�#���!192�.168.0.1�0����CAMPRYTs�O�!c�1l�����RT������ׄNAME !~�!ROBO���S_CFG 1�d� ��Auto-st�artedtFTP%�<>�� r�/A�e w����R��0//+/�#�v� ���/���/�/�/ �/?�&?8?J?\?n? �/?�?�?�?�?�?�? '9}?jO�/�O �O�O�O�O�?�O__ 0_B_eO�Ox_�_�_�_ �_�_O+O=OoQ_>o �Oboto�o�o__�o�o �o�o'o�o#L^ p���_�_�_o  �Go$�6�H�Z�l�3 ������Ə؏�}��  �2�D�V�h���� ���ԟ���
��.� ���d�v��������� Q������*�q��� ������{�ݟ��̿޿ ��ɯ&�8�J�\�n� ��Ϥ϶��������� E�W�i��}�j߱��� �߲����ߝ����� 0�S�T���x�������T( _ERR �f2
����PDU�SIZ  b�^�����>�WR�D ?qB�� � guest`�P�b�t��������!SCDMNG�RP 2gq���B�b�[$�`�K�� 	P0�1.02 8'� �  ���  � @  �
=� ����wG�*���u>G �����7�ﰀk���4�Zw ��B(Ї7��)����� r~������y�+�-�"C�l�
d-?Q��__GROU��h������	���QUPD  >ղ����TYf �����TTP_A�UTH 1i��� <!iPen'dan��,.k��!KAREL�:*,/5/G-KC�\/l/~/T VISION SET��/�/b�R"�/�/? Q#/??G?A?�?e?w?��?�?�>�CTRL� j����Eb�
�b�FFF9E�3�?@�FRS:DEFAULT:L�FANUC �Web Server:J(B�8�J��<��O�O�O�O�O_��W�R_CONFIGw k�� :O���IDL_CPU�_PCY@b�B��C�xP BH^UMI�Ni\(�|UGNR_�IO���b���`PN�PT_SIM_D�O�V�[STAL�_SCRN�V ���INTPMOD�NTOL�W�[�AR�TY�XxQ�V� �E�N� �U�\TOL_NK 1l��L� �o�o�o�o�o�o�odbMASTE�P�db�SLAVE m���uRAMCAC�HE
bO!O_�CFGLccdsUOx�o`rCYCLK�~uS@_ASG 19n��*�
 �o� ��'�9�K�]�o����������ɏۏ�k�rN�UM���
`rI�PI[wRTRY_CNY@�R��`r�Q��a��� `r�pir�o*~D�D�`PS�DT_ISOLC�  ���$J_23_DSLdN���OG�1p*{�<��<zPE�?��,��?�	߂�Q������ʯ��� ��$�`�Οؘ��PheqC�ޒPBpECMo~�UKANJI_p� �_��Z MON #q�_b�y�π�&�8�J��X"��r�;\FlŇ���CL�_L�P�$���EY�LOGGINlp�D������$L�ANGUAGE Y�F;bSD �6��LGjqs�y`a� �b�xC��G�J@~P�b�'0*_�b�;b�=MH� ;��
��(UT1:\ZϤߥ �߷���������#�L�G�Y�~�(�����LN_DISP �t*q؀�~���O�CboRDz�S�A��OGBOOK u'��������Xp�i�{��������O*3�K���F	+�r١Bs�(:s�����_BUFF 1vom?�J@ tD� B�CG��� ��!*WN` ���������/��XDCS yx�{� =����� !��E�/�/�/�/4$�IO 1y�{ ���#�0��/?? (?<?L?^?p?�?�?�? �?�?�?�? OO$O6O�HO\OlO~O�O�O�%E�PTM��dB��O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o�AoSoeo��BSEVtd����FTYP����O�o�o�otm��R�SB���V\�FL 32z�-j��e/e�w�����T�P�����b�NG�NAM�%�0$UPS��GIB���o��@�_LOADP�ROG %��%�PLACE_S�ALIDA���MAXUALRM�p�A���F�_PRB��f� ���C���{'��������Pw 2|�� ؄�	�a�
*eЃ ��X���o�����c( ���ԟ���C�.� g�R������������ ȯگ��?�*�c�u� X������������޿ ��;�M�0�q�\ϕ� xϊ��϶������%� �I�4�m�P�bߣߎ� �߲�������!��E� (�:�{�f������� ������� ��S�>� w�b����������������DBGDEF �}�u!���� _LDXDISA+���{�#MEMO_A�P%�E ?�{
 "�~����������IS�C 1~�y��� ��IS�'_������+_MSTR� �m�SCD 1�m��./� R/=/v/a/�/�/�/�/ �/�/�/??<?'?L? r?]?�?�?�?�?�?�? O�?�?8O#O\OGO�O kO�O�O�O�O�O�O�O "__F_1_j_U_g_�_ �_�_�_�_�_o�_o Bo-ofoQo�ouo�o�o �o�o�o�o,P ;t_����������:��MJ�PTCFG 1���7����[`�M_IR 1����J�@�K�̏ޏ��< ! ?�����N��K� �C�e�g�y���ɟ� ������ҟD�&�0� R���*���������ܯ 
����K�]��� ��f�p���̿j�Ŀֿ ����J�,�}Ϗϡ� 4�V��Ϫ�����߮� �F�,�>�`�b�p��� ��f�xߚ������� T�:�\��p����� �����������2� <�N�`�~��������� ����I[��� d�v���h��� �H*{��2 T����/�/�D/*/</^/�/n]�Kvc��i�  �/~[�LTARM_�"���x �"w�n��?4]�METPUw  o"���%�\�NDSP_AD�COL25� =>CM�NTS? F5MST ��-�?w��!��?�4F5POSCFzs7~>PRPMr?��9STQ01�i�4��<#�
AA5�AE QO_G=O_OaOsO�O�O �O�O�O�O!___W_ 9_K_�_o_�_�_�QF1�SING_CHK�  V?$MOD+AQ�#�i��,�.~�UDEV 	i��	MC:1lHS�IZE20�-��UT�ASK %i�%�$1234567�89 �o�e�WTRuIe��i� l��%��og�o)}��F�cYPkaz�d�S�EM_INF 1���'a`)�AT&FV0E0�2�})�qE0V�1&A3&B1&�D2&S0&C1�S0=�})ATZ���tH�)��qQ��xAY���<�����ɏۏ � ��� ��Z��~������� g�؟�������2�� ��h��-�?�����u� ��
�ůϟ@���d� K�����M���q����� ���˯<�s�M�r�%� ��QϺ��ϳ��ϣ��� &�ٿ���n߀�3Ϥ� ���߃ߍ��߹�"�	� F�X��|�/�A�S�e� ������C�0���T���e���q���*oNIwTOR�0G ?Ek�   	EX�EC1o"��2��3���4��5���`��7*��8��9����x� \��\\\ \&\2\>\J�\V\2c2o2�{2�2�2�2��2�2�2�3�c3o3�QR_�GRP_SV 1݊~{ (�Q?�������;��j�o!��"{��,m�a_DM�nn��ION_DB`�|mo!  ��0� h��+���! h��N l� }" i-ud1We�m//�/�!PL_N�AME !�e�� �!Defa�ult Pers�onality �(from FD�)<"*0RR2u �1�L68L�@P�!%`
 d �2??+?=?O?a?s? �?�?�?�?�?�?�?O O'O9OKO]OoO�O��2?�O�O�O�O�O_ _*_<_N_��<�Ox_ �_�_�_�_�_�_�_o o,o>o=,��g_xn
go�o��P�o�o�o �o�o"4FXj |������o�o ��0�B�T�f�x��� ������ҏ����� ��P�b�t������� ��Ο�����(�:��L�^�p� Fs�  GT�G��M���  �������d����ί� į����u�p���G�pX�B�{�~� k� ��������οԿ�Ϡ��7�G̛�k�	�`��zόϞ�]�:�oA<)�����ϙ� A�  	٤�"�#��)2 h�?, � �� ~;� @D�  Nу?�T�:�,!Vћ�A�/��N�Un��;��	lf�	 �xJ�Ќ�3 4 �� �<� ���� ���ґK�K ���K=*�J����J���J9�]��\�����@�t�@{S�6��(EB�n������=�N�����Il�T;f��a���������*  ´  �V �>�����T����>����ӧ�U��x`j�� ����g���j�4!��}���  {�  @.����/  �" �F�j��d��	'� �� ��I� ��  �
Ш�:��È��È=��Q;�
�[��( �5�?�n @����@���i�@�����x�;!P  'f�3�g�@2��@�W0@s�@w�@{��C��C< C���\C��C��C��^!!�@���f� ��d0�B< �	�0����&��Dzc�I���mX}�
���( �� -��������A��;��  �����?�ff!�//�� W�K/]+�8��s/�*>��<�b��	(���%P�(��ѮӼ��?����x����1�<
6b<�߈;܍�<��ê<���<G�^���#?��A���U��@�f��?f7ff?9�?&`0.��@�.r2�J<�?�\�~2N\� ���[1g��Vն?T� �?D7��5/
O�?.OO RO=OvOaO�O�O�O�O�ȟ5F���O_�O�0_�?Q_�9#_�_XG�@ G@0��G�� G}��s_�_��_�_�_oo@o+o+BL��Bh�AQo5o �o�m-�m�o���K_ o_8�o\n���|��b���#/A @|J�F���=�/ù�A� Z����A*���&��ߞ�?�ؽ�ď��菦���W�����CP�K�CH�BZׄj�y�ցz�@I�Vn�(hA� �A�LffA]��??�$�?��!��°u�æ�)��	ff��Cϼ#�
^���g\�)�2�33C�
������<������G�B����L�B�s����	�"��H�ۚG���!G��WIY�E���C�+���I۪I��5�HgMG��3E��RC��j=R�
�pI����G��fIV�=�E<YD �S�����ۯƯد� ��5� �Y�D�}�h��� ����׿¿����
� C�.�@�y�dϝψ��� ����������?�*� c�N߇�r߫ߖߨ��� �����)��M�8�]� ��n���������� ����I�4�m�X��� |������������� 3WB{fx�������(ξ����?�"��<^��N`��3�8�z����4Mgu������VwQ��4p�+4�]��>/@,/b/P/�/t,�eP2	P�.�a�o�/4�/0??;?&;RA?H?`�?l?�?�?�?  ��?�?O�?)OOMO��/�o�OnO�O�K �O�O�O�O�O __$R&_8_n_\_�_�_�_��Z  2 Fs޵�GT��V��M��B)�V�c�J�C�pc@g�,o��ISo�eo8o�o�o �\!��WɃ�o�o�o~z?���@@z��T����EA:����
 s ����������'�9�K�]���Mq �����D���$MSKCFMA�P  �� �VMqIq���ONREL  ��%���P��E�XCFENB߇
8��х��FNC���JOGOVLI�P��d��d��KE�Y߇K�T�_P�ANވf�b���RU�N;�g�SFSP�DTY� ��ӃS�IGNߏ�T1M�OT=����_C�E_GRP 1����\>OB�6O f�x��Tb���Z�ǯ~� ������!�د�W�� {���D���h�տ翞� �¿�A���e�w�^� ��RϿ��ϸ��ϡf��QZ_EDITܔ���уTCOM_C_FG 1���Xv�P�b�t�
0�_AR�C_���%*�T_MN_MODEܖ��
�UAP_C�PL���NOCH�ECK ?�� �%����1� C�U�g�y�������������	��ȋNO_WAIT_Lۗl%��NT8����zO{m�_ERR�s2����Q� ����������|� ��Բ�O���| ��BB������$���v���\T�¤ؑ��_ ��<��h?��l�%Hp����PA�RAM�򙣋�	��N8�_8� =�P345678901RdvM �������/%/+N7�W/i,���/тODRDSP���ޖ
�OFFSET_CAR����&�DIS�/�#S_Aβ�ARKܗ&�OPEN_FILE� �B�v�&֎�OPTION_IO\�n�G0�M_PRG %���%$*�?�>#3WmO0� �
!� �5���2��
r�0~'�1	 �����3������ RG�_DSBL  ģ��P|LO�!RI_ENTTOހ���C�Gp��a� UT�_SIM_DO7誂}�� V� LCT �w�"��4v��Ix��S��A_PEX����/�DRAT�� d�
��D� UP )��N^p!��C_U_2r@S:�Aq�RH�W]��$�2��L�68L@P�C
 d}/�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o $6��2�_fx� �������} U2�D�V�h�z����� ��ԏ������"� 2�pP2�X���PE��� ������ʟܟ� �� $�6�H�Z�l�~���_� q�Ưد���� �2� D�V�h�z�������¿ Կ����
��.�@�R� d�vψϚϬϾ���������߮��O'�W�i��C#�ߙ�~� ����<�<�|/���1����0&�P�F�X�j� ������$sQ���&�	`:�4�F�X���:�o{Av��������%A�  ����T�PO)P1�[�v�T}"�, �D�[0�� @D�  �����?�D�� H;�	�l�	 ��xJf ��9:]  �<w �| � ���$H(��H3k�7HSM5G�2�2G���GNɁ3�HI���$C%fp@ap@���,�Q#ã0�s@�4
*>**�9/��A�q½{=q�ª��Pd ��%�$����;$���@{ � @k@�P0�  ��0�&$�"/�P%	'� � �@"I� � � ���f=����d/v+��� � ���n �@�"�A�/'+B�$���N|@? C 'R0&4��0C|@_C��\CYC]�Ca3?E?��0�K@�
f�0�d�P�B|@�1�����!�5(z�Of+OO;O�aO��( �� -P"�!A!x�1�E�S  ����1~Qzр?�ff0���O�OfO �	_D[MA8�1_?Z>�!H�� DJ(�mUPvX��Isll�#?�՚�x���<
�6b<߈;����<�ê<�?��<�^¤�_2�AA�+��#$���?fff?�?y&`�@�.0b�J<?�\�<bN\�AI�2a
M@ to�ogX�O�o �o�o�o�o4X jU��w����_o�o�o�B��xG�@ G@0�G�� G}t�1���}������ڏŏ���BLy3B"�A��T� ?��/��I�?�#	�ϟ -���A��,�>�P��F��b�I7�OA @|����ů��¯���s�A�0��?y5�C�M��>\�?Ƀ�{�������ѹ�mWy3��οC F	�CH˿ ���������8�@I��(�hA� �AL�ffA]��?��$�?�yQӺ���u�æ�)��	ff��C��#�
�~�g\)�Pb�33C�
������<��p�G�B����L�B�s?����	�RӺ�H�ۚG��!�G��WIY�E���C�+��нI۪I�5��HgMG��3E��RC�j�=�
�pI����G��fIV=�E<YDf� Կu�`ߙ߄ߖ��ߺ� ������;�&�K�q� \���������� ����7�"�[�F��j� ��������������! E0iTf�� �����A ,eP�t��� ��/�+//O/:/ s/^/�/�/�/�/�/�/ �/? ?9?$?6?o?Z?@�?~?�?�?�?�>(p�g���o�R��E�5��OOa��3�8�8OJOa�4�MgudOvOa��V�wQ�O�O4p�+4�]�M�I�O�O� __D_2\��P�RPv^�����_�?�_�_�_�_�[R�_o?o�*oOouo`o  �@� xo�o�o�o�o�o�_`��>,bP{h�r������� ��,��P�>�t���  2 Fs_��GT����M�a�B���!��C�.�@%����� �2�D�U�����������ǟa�?���@U@Κl�a�a��o�a�p�
  Ο1�C�U�g�y����� ����ӯ���	��r��� ��`K�D���$PARAM�_MENU ?��E� � MNUT�OOLNUM[1-]]�v�FX�]���AWEPC�R��.$INCH�_RATE��S�HELL_CFG�.$JOB_BA�S�� WVW�PR.$CENTER_RIϲ��ִ�AZIMUTH �OPTB��ִE�LEVATION� TC��ִDW���TYPE SN���ARCLINK�_ATڰSTAT�US��7�__VA�LU����LEP>�.$WP_}��� gU��|ώϠ������π�����0�Y�T�S�SREL_ID � �E�Q�h�US�E_PROG �%c�%Uߺ�i�CC�RTxԐQk���_H�OST !c�!�����T�P��+�����-�g���_TIMEOU��g�	�~T�GDEBUGx��c�i�GINP_FOLMSK���T`l����PG>�  ��n���CH���+�
a�l�T�N߄��� ����������= 8J\����� ���"4] Xj|��������/5/��WOR�D ?	c�
 �	RSe	PyNH��2MAI1�fp#SU �|#TEN�>�3STYL�s �COL
e1(�/1�T�RACECTL �1��Em� �tP�P�'DT �Q��E0� D� � fS��r+6�5;K?]? o?�?�?�?�?�?�?�? �?O#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �_�_�_�_�_	oo-o ?oQocouo�o�o�o�o �o�o�o);M _q������ ���%�7�I�[�m� �������Ǐُ�����!�3�E�W��&LE�1�z����#  ���&_UP ��;<�����ñ ��� �� ��$;�ޟ��60�  ���)_DEFSPD� �c�2�� � �T�IN��T�RL ���;�8���B�PE_CON�FI����'�t��!<,LID������	��GRP �1��) l�V�@�j��h�s�!A�
D��� D@� C�o� @��^� �d���)������ྠ"�����C� ´|�^�G�B�����p����������!>��>�,���7�I��3� =49X=H�9Nχ�JτϽϨ� ����f���)���9�_�J�  Dz�Ӎ�� 
tߵ�d�������� ��3��W�B�{�f�x�@����������)��
V7.10b�eta1Ӗ �A���6��!���3�?!G�>¿�\=y�#2�{�33A!��@����2��8wA���@� A�"�@�#�B� �����������#Ap�"�����dd��$�?����@, �� �Ay��33@���#� Ҿ��/�xߋ���ǡ�KNOW_M  �
���SV ]��*�%�� ��������#��"!�ãMʣ��-���	ٕ (���ڔ@7X�#�{�3�@{����������MRʣ��-�$��`����@/R+��STʡ�1 1�98 4�
Carga_7Too}?�'/���#Pieza ����/�'��ø��/ �/
??.?@?R?d?�? �?�?�?�?�?O�?O@KO*O<O�OW�p'2{,�e4cO  �<�O�Ow 3�O�O�O�O�p'4�O__+_p'5 H_Z_l_~_p'6�_�_�_�_p'7�_ oo$o�p'8AoSoeowop'M�ADw� ���EO�VLD  ����*}p$PARNUM  ~+s��/�T_SCH�i ���
}wFq�yē�uU�PDFuY���E_CMP_Ow�Ҡ9��'���tER_CHK���ڒ!�
���RS ]��_M�O�`o���_k��E__RES_Gz ���
��J���� ��D� 7�I�h�m�������@�ٟ�o���@Ɍُ ����@(�G�L���GP g��������P��ůʯ ���P��	���@`$� C�H����`c��������V 1�ʅ��e�@]s8��THR�_INR ' dz��d��MASSϛ Z�MN�5�M�ON_QUEUE� �ʅf2�� U��N�UH�NE�nȅ�END�������EXE�Ϥ��pBE����υ�OPTIO��Ǳ���PROGR�AM %h�%�����l��TASK�_I�d��OCFG� �h�\ߏ�D�ATAR����'2p���"�4�F� ��j�|����]�����������INFOR���w�y���e�w� �������������� +=Oas������(�4���� ����ѥpK_��Ѵ��T�G��2�� X,		�R�=���d�'�@�u@}$;�`�||�
_EDIT �������WERFL���m#�RGADJ �^�A�  +%?�!�8$
�&���ʅO��,��<|n@T�%�o�/(�M#f�2�Y'�	H��l��f!?#��8A���t$6�*0/2 **�:&2n@?+3G=ʅ�`2[5��1e9΁ �/nB�?S=�=c?u?�? �?�?%O�?�?OOO �O;OMO{OqO�O�O�O �O�O�O�Oi__%_S_ I_[_�__�_�_�_�_ Ao�_�_+o!o3o�oWo io�o�o�o�o�o �o�/Aoew ������]�� �G�=�O�ɏs����� ����5�ߏ���'� ��K�]���������� ɟ�����y�#�5�c� Y�k�寏���ϯůׯ�	��p�l ^����� 9��3��濁�
���I'PREF ��Y*l l 
%IOORITY���!MPDSP�*�"�w�UTz��#&OD�UCTw�����&OG� _TG��|����TOEN�T 1�� (�!AF_INE���3�j'!tc�p>�f�!ud�Uߎ�!icmX}ߥ.��XYR#��;�l!)� 31���l ���-��� Y�@�}�d�v����� �������1��U�g�	*��R#�Y)�"�/�����l#>��F"1�B37/=<��l$��(��.A{",  �O�Wi{�%���8��@�R�	"!PORT_NUM���l �!_C?ARTREP���;SKSTA�� �LGS0�����{#l Un?othing�s���&�7TEMPG ��ɣ.�[�_a_seiban�/�/</'/`/ K/�/o/�/�/�/�/�/ ?�/&??J?5?n?Y? ~?�?�?�?�?�?�?O �?4OO1OjOUO�OyO �O�O�O�O�O_�O0_ _T_?_x_c_�_�_�_��_�_�_�VERS�I����'` disable����SAVE ����	2670H�771���_�o!`���o�o�߻o 	�hH��0�{��e% N`r�$�=|�o����Gb_�� 1�
��p`�J����� ���1�URGE_�ENB������W�FL�DO�Ƥ�W�,�m���
WRUP�_DELAY ��`�R_HOT %U������~��R_NORMAL�̈��܏1� �SEM�I�6�u�/�QSKKIP�sƺ�sx�_ ���_ޟ��ŝ�3� !�W�i�{�A������� կ�������A�S� e�+�u�������ѿ� ������=�O�a�'� ��sϩϻ��ϓ�������'�9�K�υ�$R�BTIFn�
RC_VTMOU�ջ�i�DCR�sȾ�� �ё6���CB}�C�jP>�Cg>��9L�&ŝ���e�cw����R�E���ş��� <
6b<�߈;܍�>u�.�>*��<ȃ��'�� �z�� S����������	���-�?�Q�c�u��RD�IO_TYPE � �}k��EFP�OS1 1�Oi� x�o
�h�! E�oi�(�� ^���/A� �(�t�H�l ���+/�O/�s/ /�/�/D/V/�/�/�/ ?�/9?�/]?�/Z?�? .?�?R?�?v?�?O�?��?�?YODO}O��OS/2 1ʮ���4O�nO�OjO_�O��3 1˨O�O�O_�_o_|�_&_S4 1�=_�O_a_�_oo=o�_S5 1��_�_�_0o�o�o�oPoS6 1�goyo�o�oC.g>�oS7 1��o� Z���zS8 1Б���m��X����SMASK 1ў� ��ЏچN��XNO��͆�<���MOTEp������4�_CFG ��;������PL_�RANG7�s�u�O�WER ��������SM_DRY�PRG %��%�8�����TART �Ԡ��UME_�PRO��ϟJ���_�EXEC_ENB�  `�{�GSP�D#�e�m���|�TD�B����RM����I�A_OPTION�ּ�}�/�MT_"��T��9���T����c�C������[�m����\�i�O�BOT_ISOL�C��j�g���N�AME ���9���OB_ORD_NUM ?�����H77�1  ��B�@�B���Bʆ�B��PC�_TIME��w�x�i�S232T�1����̱LTEA�CH PENDA1N��P��X�7��"@Mainte�nance CoKns���ϔ�"���DNo Use X����C�U�g�yߋ����NPO����������CH_Lf&��/���	�~��!UD1:3�z��R��VAIL#�����/�SR + ����o����R_INTVAL�������ꮅ�V�_DATA_GR�P 2�����2�D��P��1��U�@� ��x���p��������� ������ H6l Z�~����� �2 VDfh z������/ 
/,/R/@/v/d/�/�/ �/�/�/�/�/??<? *?`?N?�?r?�?�?�? �?�?O�?&OO6O8O JO�OnO�O�O�O�O�O��O�O"__F_/��$�SAF_DO_PULS��0���2�pQN`PCAN������SC�����(����G��K����PR������ J� �_
oo.o@oRo�_vo��o�o�o�o�o��J��kb2�dڍd�d�qF�s�� @�n�@Rdv~(y� ���t�_ @�T������~��T D��� -�?�Q�c�u������� ��Ϗ����)�;��M��߱�:u��������o���¯;�o����p����
�t���Dia�la�Q��  � �Ϻ�QlaR� �Q;�M�_�q������� ��˯ݯ���%�7� I�[�m��������ǿ ٿ����!�3�E�W� i�{ύϟϱ���������ߕ��;4�F�X� j�|ߎߠ߲�����e ����&�8�J�\�n� ������r0�� �(�������+�=� O�a�s����������� ����'9K] o������� �#5GYk} �������/ /1/C/U/g/y/�ߝ/ �/�/�/�/�/	??-? ������kbm??�?�? �?�?�?�?�?O!O3O AITOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�_�_�_�_�_�_@�_oo(o:o��c� �Eo�o�o�o�o�o�o �o $6HZl~��Jjoo��.����-��_��	123456�78�h!BO!ܺ[4��m`��V�h�z������� ԏ��no�!�3� E�W�i�{�������ß ՟�����/�@��� c�u���������ϯ� ���)�;�M�_�q� ��B�T���˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����Ϙ����!� 3�E�W�i�{ߍߟ߱� ����������/��� S�e�w������� ������+�=�O�a� s���D���������� '9K]o� �������� #5GYk}�� �����//1/ �U/g/y/�/�/�/�/ �/�/�/	??-???Q?c?u?�?NcG��?�?�K/�?�?O �C�z  BpKj  W �]h2abG��} Lh
]G�/  	�Nb2�?�O��O�O�O�K>�9DFo�<�wO_._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro _�o�o�o�o�o�o &8J\n�� ������I.B��1kACB<-���$SCR_GRP� 1��8�� � � ��.A >E	 b��j�{�t��1���,G�������܏M�,M@قD�W�N����ً�L	M-1�0iA/7L 1�23456789�0m@P� 8m@cMTW�_�.C
Z�����\�]KSB��_ j�.FY���Y��Cف�Ax�����	SJ�"��4�F�X�.D��#H�j��n�Y��������ǯٯ���o.A �����A��3�p���B�'@ƌ�������9A8@��  @.@ʵD���?�@򵆲H'@��ݺ��F@ F�`-�5�,�Y�D�}� hύϳϞ�������~��ʱ��&��#�5�G�B�U��ϛ߆߿ߪ��� ������=�(�a�L� ���O���ŏ����>G�_@��
�.B�ʱ6G�.��Ȱ��@ʰ4J�'@�`�Z���0���?��.DA�����$�����A��.AA ������B�N`/ (�  ����}�����.F9�EL_DEFAULT  Ô���.@~HOTSTR&���:MIPOWE?RFL  E2�`WFDO'� tRVENT �1���s�Q� L!DUM_�EIP,H�j!AF_INE&<�.D!FT�.��>/!��c/ ��-/�/!RPC�_MAIN�/m(�8y/�/�#VIS�/l)y��/"?!TP0�PU?�d?n?!�
PMON_PR'OXYo?�e]?�?�52�?�f�?O!RDM_SRVOr�g�?RO!R��dnO�hAO�O!
� �M�?�i�O�O!?RLSYNC�O���8�O6_!RO�S�]\�4%_�_!�
CE70MTCO�M�_�kq_�_!	��RCONS�_�l�_o!�RWAS�RC!O�m	ofo!��RUSBgo�n Uo�oQ/�oC�o�o�o $�oHl3��RVICE_KL� ?%� (%�SVCPRG1�����u2���p3����p4/�4��p5�W�\��p6����p7@�����p{���|9�����tiO$��q�L� �q�t��q!����qI� ğ�qq���q����q ��<��q�d��q��� �q:����qb�ܯ�q�� ��q��,��qڟT��q �|��q*����qR�̿ �qz����q����ʯ ��r�p��pgϬ��q ���Ͽ�������@� +�d�v�aߚ߅߾ߩ� ��������<�'�`� K��o��������� ���&��J�5�n�Y� �������������� ��4F1jU�y ������0��z_DEV ~��MC:o��4��JGR�P 2�o��p�bx 	� 
 ,�8�o �� /��6//Z/ A/~/�/w/�/�/�/�/ �/?�/2?D?�h?? �?�?�?�?�?�?�?�? OO@O'O9OvO]O�O �O�O�O�O�OK?�O*_ �ON_5_r_�_k_�_�_ �_�_�_o�_&o8oo \oCo�ogoyo�o_�o �o�o�o4-j Q�u����� ���B�)�f�x��o ��S���ҏ����ݏ� ,��P�7�t�[�m��� ��Ο�����(�� �^����i������� ܯï ����6��Z� l�S���w�������� A�� ��D�+�h�O� aϞυ��ϩ������� ��@�R�9�v�]ߚ� ����߇������*� �N�`�G��k��� ���������&�8�� \���Q���I������� ������4F-j Q���������id �i	 U@yd����)%���q����!�%/,'/ L/:/p/^/�/�)��/ 
)�/�/�/??(?*? <?r?�/�?�/b?�?�? �?�?OO$Oz?�?qO �?JO�O�O�O�O�O�O _RO7_vO _j_�Oz_ �_�_�_�_�_*_oN_ �_Bo0ofoTovo�o�o �oo�o&o�o> ,bPr��o��o �����:�(�^� �����N�p�J���� ܏� �6�x�]���&� ��~��������؟� P�5�t���h�V���z� �������(��L�֯ @�.�d�R���v���� ��$�����<�*� `�Nτ�ƿ���t��� p�����8�&�\ߞ� ����L߶ߤ������� ���4�v�[��$�� |����������N� 3�r���f�T���x��� ������������� ,bP�t���� ��(^ L����r��  /�//$/Z/��/ �J/�/�/�/�/�/�/ ?b/�/Y?�/2?�?z? �?�?�?�?�?:?O^? �?RO�?bO�OvO�O�O �OO�O6O�O*__N_ <_^_�_r_�_�O�__ �_o�_&ooJo8oZo �o�_�o�_po�o�o�o �o"F�om6 X2������ `E���x�f����� ��ҏ����8��\�� P�>�t�b�������Ο ���4���(��L�:� p�^���֟��ͯ���  ��$��H�6�l��� ��ү\�ƿX�ֿ���  ��Dφ�kϪ�4Ϟ� ���ϰ��������^� C߂��v�dߚ߈߾� ������6��Z���N� <�r�`�������� �������J�8�n� \������������� ����F4j��� ��Z������ B�i�2�� �����JpA/ �/t/b/�/�/�/�/ �/"/?F/�/:?�/J? p?^?�?�?�?�/�?? �?O O6O$OFOlOZO �O�?�O�?�O�O�O_ �O2_ _B_h_�O�_�O X_�_�_�_�_
o�_.o p_Uogoo@oo�o�o �o�o�oHo-lo�o `Npr����  �D�8�&�\�J� l�n������ݏ��� ���4�"�X�F�h��� 䏵�􏎟�֟��� 0��T���{���D��� @����ү���,�n� S������t������� �ο�F�+�j���^� Lς�pϦϔ϶���� �B���6�$�Z�H�~� lߢ������ߒߴߎ� ��2� �V�D�z�ߡ� ��j�����������.� �R���y���B����� ����������*l�Q ���r���� �2X)h\J �n���
�. �"/�2/X/F/|/j/ �/��//�/�/�/? ?.?T?B?x?�/�?�/ h?�?�?�?�?OO*O PO�?wO�?@O�O�O�O �O�O�O_XO=_O__ (__p_�_�_�_�_�_ 0_oT_�_Ho6oXoZo lo�o�o�oo�o,o�o  D2TVh� �o�����
� @�.�P������v� Џ������<�~� c���,���(���̟�� �ޟ�V�;�z��n� \�������ȯ���.� �R�ܯF�4�j�X��� |���Ŀ��*���� �B�0�f�Tϊ�̿�� ��zϜ�v�����>� ,�bߤω���R߼ߪ� ��������:�|�a� ��*��������� ���T�9�x��l�Z� ��~��������@� P���D2hV�z �����
� @.dR���� x��/�/</*/ `/��/�P/�/�/�/ �/?�/?8?z/_?�/ (?�?�?�?�?�?�?�? @?%O7O�?O�?XO�O |O�O�O�OO�O<O�O 0__@_B_T_�_x_�_ �O�__�_o�_,oo <o>oPo�o�_�o�_vo �o�o�o(8�o �o��o^����  ��$�fK���~� �������؏Ə��>� #�b��V�D�z�h��� ����ԟ���:�ğ.� �R�@�v�d������ ӯ������*��N� <�r�������b���^� ̿��&��Jό�q� ��:Ϥϒϴ϶����� ��"�d�I߈��|�j� �ߎ߲߰�����<�!� `���T�B�x�f��� ���(���8���,�� P�>�t�b�������� ������(L: p�����`��� ��$H�o� 8�������  /bG/�/z/h/�/ �/�/�/�/(/??�/ �/�/@?v?d?�?�?�?� ?�?$?'1�$SE�RV_MAIL � .5$@�
HO�UTPUTH�
HRV 2��6  '@ (�1�?�ODTOP1�0 2�ZI d *?�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����5�E�YPE:L(EFZN_CFG �5�'C'4IB�xG�RP 2��w�q ,B   A?�~'1D;� B@���  B4'3�RB21�FHELL�r�5�vm@nO�����;%RSR����ʏ��'�� K�6�o�Z�l�����ɟ����؟�#�5��  ��5�c�u�,C��� '0}���(��'8K�2'0d����|�j�HK 1�x� ���$��H� q�l�~�������ƿؿ ���� �I�D�V�h�~d�OMM �x����i�FTOV_E�NBDbA�u��OW_REG_UI���BIMIOFWD�L����B��WAIT��٩IE8�4@r��aD2�TIM��7��l�VA@C�>�_UNIT�ã�v�yLC��TRY����u@MON_�ALIAS ?e��i@he�?'�9� K�]�%:������ o�������0���T� f�x�����G������� ����,>Pb s����y� (:�^p�� �Q��� //� 6/H/Z/l//�/�/�/ �/�/�/�/? ?2?D? �/h?z?�?�?�?[?�? �?�?
O�?O@OROdO vO!O�O�O�O�O�O�O __*_<_N_�Or_�_ �_�_�_e_�_�_oo �_8oJo\ono�o+o�o �o�o�o�o�o"4 FX|���] ������B�T� f�x���5�����ҏ� �����,�>�P�b�� ��������g����� �(�ӟL�^�p����� ?���ʯܯ� ���$� 6�H�Z��k������� ƿq����� �2�ݿ V�h�zόϞ�I����� ����
ߵ�.�@�R�d� ߈ߚ߬߾���{������*�<����$S�MON_DEFP�ROG &����f� �&*SYSTE�M*C���R �S�RECALL �?}f� ( ��}2xcopy �fr:\*.* �virt:\tm�pback��=>�192.168.�56.1:928�4 ������.�}3��a�������������>�7��s:o�rderfil.datP�b�x�	�-}.��mdb:M���4 ����� 9���T���w, ?���u������ ��Xs//(/;M ���/�/�/�L^ � ??$?7I�/m ~?�?�?��P/��? O O3/E/�?i/zO�O �O�/�/V?�/�O
__ �OA?�Oe?�O�_�_�_ �?�?ZO�Ooo*o=O �_aO�_�o�o�o�ON_ `_�O&9_�o�o o_����_�_Ro�_ ��"�5oGo�ko|� �����o�oX�o��� �1Cԏg.����� /���\�w���,� ?�ڟc����������� P�]����(�;�̯ ޯq���������˟T� � ��$�7�I��m� ~ϐϢϵ�ǯZ���� � �3�E���i�zߌ� �߱�ÿտc߮�
�� ��A���e��߈��� ��R�_�u���*�=߀����s߄�������6�B�:pick_e�ntrada.tpP�emp\�w��+��4��index���������� }5��lace N`��(���sali���.� ������[�u// +/>��b���/�/�/���$SNPX_�ASG 2������!�o  0�%��/��/  ?��&PA�RAM ��%��! �	�+Pʴ��I4��� OFT_KB_?CFG  ��%��#OPIN_SI�M  �+D2��?�?�?�3� RVN�ORDY_DO � N5v5�2QS�TP_DSB�>�D2"O�+SR �>�) � &H:eO���&TOP_O�N_ERR�?�FP_TN �%�@��C�BRIN�G_PRM�O�2V�CNT_GP 2���%F1� x 	 O_�_@_+_d_�'�VD�@RP 1�9G0UQ�1G_�_�_ �_�_�_ooo/oAo Soeowo�o�o�o�o�o �o�o+=Oa s������� ��'�9�`�]�o��� ������ɏۏ���&� #�5�G�Y�k�}����� ��ş������1� C�U�g�y��������� ӯ���	��-�?�Q� x�u���������Ͽ� ���>�;�M�_�q� �ϕϧϹ������� �%�7�I�[�m�ߑ� �������������!� 3�E�W�i����� ����������/�V� S�e�w����������� ����+=Oa�s}RPRG_CO7UNTk6�B�	'ENB�O�M�m4��_UPD 1�>HKT  
�� -?hcu�� �����//@/ ;/M/_/�/�/�/�/�/ �/�/�/??%?7?`? [?m??�?�?�?�?�? �?�?O8O3OEOWO�O {O�O�O�O�O�O�O_ __/_X_S_e_w_�_ �_�_�_�_�_�_o0o +o=oOoxoso�o�o�o �o�o�o'P K]o����� ���(�#�5�G�p��k�}�������ŏ�_INFO 1�	�  �� �,���P�;�����?�?0*?��V�=��B����������˘=K%��¤؏³����YSDEBUG�� 
�׀d�	��S�P_PASS��B?̛LOG ��	  r׀׈�  ���ׁUD1:\x�����_MPC���	z���	5��� �	Z�SAV ����B�!�9�ׅ�@�SV��TEM_TIME 1��] 0� ���ά�L��SKMEOM  	�!�  ׂ%M������ׄ� @׀� �(ׂ�ׁ"�e��� A��ĲϹ�0�׃HʰׁB�nπ�ȒϤ��^��� � 	W��κp����)� ;�M�_�q߃ߕߧ߹������L���%�7� I�[�m������� �������!�3�E�W��i��T1SVGU�NS�'���~�ASK_OPT�ION� 	�����_DIې���B�C2_GRP 2��	�+���ׁ@��  C�׉A���*�*׀V9.�0055 C1/�31/2017 �A w�11M����_ACC_T���X-$tLEN1  �}2�EL_RA���� $��W_AX[IS�F1tI�=2�MOVE�����ERTIA �  	$D�T�ORQUEs�D�E��LACEMCNT�t ��V� �MAXAAT�CVHiTRQxh�STAT1��J_���M�� J_MOD��$D� T��2�P��!� JK&VKЈ1!�1!3##J0lF$5#JJ=#JJE#AAL5#k =#k e&e4f%5��N1�М [E�L� _N�UM�׀oCFG�w ` $GoROUPDSK��B_CONFLI�C�� REQUIRED����p�7$T2 -1q �6oSG��w �\ $ENAB�L�$APPR�#0CL�
$OP�ENj8CLOSEy:S_M��� �9�
oPARA� o �b0MCDx���4_MGN�3C��AV�9�C�7�BRK�9NOLD��6SHORTMO�_LI�!#GM�5J,@DPm$#=##E#�#�##�##6ZE7:ZE8���oM4�  2����G��CPATH �G�A�C�A��C�020]� CNTj0A^2�#Gk2�1INsUCh� �3PC�UM<X�Y� 0�CQYP_�E� ^Z� ^ZE ^PP�AYLOAGJ2�L_UPR_AN1�SLW�[�Q�Y�Q��5R_F2LSHR��TLO�T2Q�W�@S�W@SACRL_��0U#`,W�T�HV�Am3$H�2QbF�LEXm3o J���w PW2B_�� �!� M_FT�M��d�RESECRVjQ�g�jE!�A}Js :� ��g�d�����F1�aHu\w�@��+�rE5 GYk}���� c�����$pp�����
/�a*T��a�X <pi�%�t�x(%1�
� 4/F/X/j n%w%e%�%��/�/�/�)�BJ�$ � �/�/?�UPDATuv1�CEL�p+�F�&8JP�-0JE
@CTR,,QpqTN�pFC�7HAND_VB�r�maOPL5 $�ՀF2�6�3]�CO�MP_SW�'�6	?� $$M�P�9R�3��	A��p��B&"�A_�R�6D<��=UA�<A�<AKAKTJ��;D�<DKDK�P�@GR�7�ST��7�	I�NHDY �Ph0�6+�R��Pu �W �a�W�Q�W'��"p�EPbEkEtE}E�E�E�E�B�"JL5
 ��d�B �q�Ŝ1���ASYMUh`���V	#�"]�Q'__SH�"1WKT5M7Ի� U_g_y_�_�SJ�\U@�Z�����Y�t_VI➣�3$�V_UCNI�S8�Z��QJ % Q��Q��\U�eb�� m�'iU@6oHo����^dfc�BO0HR_T\2�����a1DI@ƃO&��B�V�#��Y�I<�A�1@SS�vpa�a��p�S�l`�p	�  �� ̡ME�qЮ�|���c�T�PT@��ؐ�@��� �Y0��Щ����T���!� $DUMMY}1b�$PS_sp�RF5p! $��n�0FLA� YPŃ���$GLB_T��4��`1�@�pt�B� XW07M1�ST�q-0SBR�PM21_Vg�T�$SV_ER�PO���z�CLN zA��pOV��GL�E�W�! 4� ��+$Y/rZ/rW� ��QȣA}�<R뒿U.� ՀN� ���$GI��}$�� � �� �!� L� ��}$Fz��E NEAR�p�NzsFg�pTAN9Czr��JOG)pK@� � $JOgINT��p���MSET�!  "EM�q�S�|��!� qp�U�q?�-0LOC�K_FO�Pӡ"�B�GLVw�GL(T?EST_XMm0�'EMP�g�5"L��$U�`��2,1�[!&"Ϡ [!�|CE� )|  �$KAR'�M(�T�PDRA� �$�VcEC�`�&�IU[!�{CHE TOOiL<s�#V;tRE� 'IS3�e�"6��pp�ACH�P�!O�P����29��� I�]2  @$RAIL_BOXE��� ROBO,$?���HOWWAR�YaK1��1ROLM q5ב4�2�90@p�@O_F�! !١� 	1�A�٠R� O�b�4p���0آ�OU��bW%��M�'��/$PIP-&NÀ�"�92	1�p[!�0�`CORDED P�1���Oc�  D 3 OB�Q� �nG]A��2 ]B��S�S;YS]AADRR����TCH� � ,ՀEN�aA
!_�D��ԣ��VWVA� Ǥ � ��PR�EV_RTt�$�EDITVVSHWR�f.P�r�%�D���aETq?$HEAD����4_P��SKE����CPSPDvVJM%Pz@L��`R�p>��e@~a�FI6 SR�C��NE� S���OTICK<sF�M��x�SHN\� @g@�Q�~Q_GqPf06�`STY�B1LON�W	b��_ t 

PG�ES%$�A=f SH�!$G����P�rP)�fSQU� x/u �TERC����R�TS� r �À����!b5�O���2pIZ!4��PRO@�+r�Q�0PU�;u_�DOl�@XS�KN�AXIZp�3`!UR ��sS�R0�P�Fdá!�_� �BET�rQP
"v@�Y`F�2Z`A����*3�$3j��SR��l�`�K���� �(�"��-��;�� K�\�m�\�}�\���n� ����n����������C���ߘߪ߼�0�SSC6    �h� DS`�!��S�PM���AT{�#��<q�P�R��ADDR�ES�#BPSHIyF�R _2CHR���AIU ڑ�TU�U I� !�COUSTO�t١V�IA�"�B(��s��=
5*
h<�HtN^ # \�PH�Y`*��a�g�C���b�r�9�F�g��TXS�CREE_B$�uaTINA�&��2�p�0Q_����% T�Q� r�A��q �hq�Bhr�PRROV���@pP ��tv�1UE�T& ����A S��ARSM<�P^wUNEX�`�q��S_���@Ӂ�����@ӜqC�m��o 2%��UE���'G�Զ+pGMTJ��Ls�wq� O�7/BBL_0W��^ �( �Y`1�O�=�LE̒H�Q0 �G��RIGHQ�BRD<�CKGR��y��TEX�pz�u�WIDTH3;Pr,1��!��UI�0E9Y��]) d� �P��=b90'qBAC�K;a/r�ū��F�OFA��LABF�?�(��I0�$UARW1,�R ����H'�� * 8��_^QڒOҎ�R� �$3�7���`<�Oӑ^ +�`�r�U]���R
"|1LUM��v��GERVA�@��Pkj��,���pGE0�hR�p�)gPLP���rE�`M�)�lQ�Pm��0�5�6�7�8���b��&pk�{���1�S��+��USR�- <�P��U�sFO��PRI�q�m#0����TRIP>51m�UN.�?�.~`.�`uc1_u��R"�p�` /�Jҹ�*qG f`T0�0;�ۑE�OS��Z�AR�p-�1��!]0�@����dO�S!U��]1��������e1�OFF+ ^ 2b z��O  10� ���"1� GU�AP�!�=8�G��SUqBb� �SRT����t3b��0
sOR�0�RAU��T��	�G�VC>�84�� /2^A�c b$��a3�C�0��DRIVv�q_�V`2P�D��MY_UBY���`f@��e9��`ҠLQo�!~P_Sz@jt �A{BMD�$�PDEY�CEX�E�&�.�p_MU�PXD����US�Q� ��� Ѡ��b���9��aG̀P�ACIN�Q�`RG Mp%#"��#"��#"����REd�Б�!�2��#"�05 �0TARG)P>�h ��Rq�06����iqd��m	�XqRE��SW _A!�$�)pO��AԐ�#��E��UL`1�V�&HKQb7`�*`�`�� �%3EA�P/7WORQ��%�0l"�MRCV�8 ����O]`MQ�C?�	pl2��e#l2REF� �6u6`1� ���s� �� q:�1�:�1�;�5u6?�_RC0;HI;��S ���5�a@b��l"�9 �.b�����`��:�`OUg`"f�� 4~%<�2�R�$��}�*p�P6蛓<��RK{pSUL6?�7��COe�f�8��@JS
�SXQ@V~�V��S�@Lz�9U�9U~�EW���|��T:| +����qՠ ��CACH5cLO�1�T�Q��Y�q���cC_LIM-I͓FR�XTt��VNVK$HOQ�mb�POCOMM�m�O[��gH��уDd�VPHb"�@Kb_vUdZ �Ph�PPhWA�UMP�ujFAI�PG!4�PAD�i�IMR1E�D�bZgGPs�����ASYNBU=F�VRTD�etlZa��OLՐD_���uW��P�ETU��PQ� �eECCUU(VEM? �Ugr�WVIRC�au�c|l�q_DELAZ#��8��kAGyR��XYZ�����W�!�s���pT� ������;����LAS���J�pQc�G�a{�<��QS�`�VN<�m��VLEXEwU=��������^cFL2v�I��cFI!p��@~��"3.�r��
t">��d�\D���\bH�ORD��������B5�?Š��T����XO������VSF��U�@ a Ǡ�Q�URR36j SM�A�2��J�����a��B�$�N�LINl��m��W�0XSK1���CJ�%�F@K��H���HOLсl���XVR
�D�	�T�_OVRт �ZABCzEz"�׃���1ZD 
�F�D/BGLVOcL5�}��ZMPCFz�GJ�k�(�}�DLN�� 
j��{�H ���a/0��C�MCM COcCAgRT_���$P_��? $JݣפD@a����s���s���"UX�q��UXE�'��q����J��0�B�0�R���ZA��I }�\��}�Y���D4� JJ�R�`���pHEk���%� �������mDK � 1��18��s�EAK�7@K_�SHIP�Vp��RVBypFv�2#��C?� آ͡�D2��>���B�If�5eDv�TRA�CEa�V�q~�S�PHER��L �,�@��п��$�TBCs� ��������  `�� �����`���	 �\�G߀�kߤߏ��� ��������"��F�1� j�U��y������� �����0��@�f�Q�����{���|����� j���%I4m���ő��a��� ���'79 K�o����� ��#//G/5/k/Y/ �/}/�/�/�/�/�(�� �/?-???Q?�/u?c? �?�?�?�?�?�?�?O O;O)O_OMOoOqO�O �O�O�O�O_�O%__ 5_[_I__m_�_�_�_ �_�_�_�_!ooEo�/ ]ooo�o�o�o/o�o�o �o�o/AS!w e������� ��=�+�a�O���s� ������ߏ͏��'� �7�9�K���o���[o ��ϟ������5�#� E�k�Y���������ׯ ů�����/�1�C� y�g����������ӿ ���	�?�-�c�Qχ� uϗϙϫ�����߻� �/�M�_�q��ϕ߃� ���߹�������7� %�[�I��m���� ��������!��E�3� U�{�i����������� ������A/e� }����O�� +OasA� �������/ 9/'/]/K/�/o/�/�/ �/�/�/�/�/#??G? 5?W?Y?k?�?�?�?{ �?�?OO1O�?UOCO eO�OyO�O�O�O�O�O �O_	_?_-_O_Q_c_ �_�_�_�_�_�_o�_ o;o)o_oMo�oqo�o �o�o�o�o�o%�? =Om���������v-��$�TBCSG_GR�P 2�u��  �-� 
 ?�  X� j�T���x�������菀ҏ��1�8��G�_d, �M�?-�	 HCA�����i��CS��B�P�����]�>'��ͱ�u�Г�۝;B��333����Bl{����#�Aʐ�fffA��5��C�#�%��s�?�����N�~�Y���A@-��ӧš����@Ư P��4����_�|�G��Y���Ŀӻ�����	�V3.00P�	Omt7���*���,��ݶY��@Wff-� -�H��� U�'�V�  ����'ϖϟ�1�+J28�?��ϫȿCFG �ueI� L������9k�*��*�P� ^��^߄�oߨߓ��� ����������J�5� n�Y��}������� �����4��X�C�|� g�y����������� P�jp);��nY ~������ "4FjU�y ��-������ /C/1/g/U/�/y/�/ �/�/�/�/	?�/-?? Q???a?c?u?�?�?�? �?�?�?OO'OMO;O qO_O�O�Og�O�O{O �O__7_%_[_I__ m_�_�_�_�_�_�_�_ �_3o!oWoio{o�oGo �o�o�o�o�o�o�o/ SAwe��� ������=�+� M�O�a���������ߏ ͏���9��OQ�c� u����������ɟ�� �#��G�Y�k�}�;� ����ů��կ���� ٯ/�U�C�y�g����� ����ѿӿ��	�?� -�c�Qχ�uϗϽϫ� �������)��9�;� M߃�qߧߕ����߇� �������I�7�m�[� ����������� ���E�3�i�W����� ����}������� A/eS�w�� ����+O =sa����� ��//%/'/9/o/ �߇/�/�/U/�/�/�/ ?�/5?#?Y?G?}?�? �?�?q?�?�?�?�?O 1OCOUOO!O�OyO�O �O�O�O�O�O_-__ Q_?_u_c_�_�_�_�_ �_�_�_oo;o)o_o Mooo�o�o�o�o�o�o �/+=�/�o m������� !�3�E���{�i��� ��ÏՏ������� -�/�A�w�e������� ���џ���=�+� a�O���s�������߯ ͯ��'��K�9�[� ��o���QϿΉ� �����G�5�k�YϏ� }ϳ������ϧ���� ��1�g�yߋߝ�W� �߯�����	����� -�c�Q��u����� �������)��M�;� q�_������������� ��7I�as �/������ �3!Wi{�K�������  9 ## #&7/�#"�$TBJOP_GRP 2���  �?�#&	O"V#
v],���� ן� =r% � ȱ � �� ��#$ @ n"	� �CA��&�?�SC��_#%n!��"G��"k���/;=�C�S�?��?��-0,0CR  B4��'F?Q7�/�/?33�3�2Y-0�?�:;���v'2�1�041*�90�=?�?90��7C�  D�!�,� �BL��O%K:��Z�Bl  @pzI@�� s33C�1y �?nO  AЁG�2qG�&0A0E�O�J�;���A?�f�f@\@�1C�a0z8qO�O�@���U�O��$fff7R0_B^;7xCsQ?ٽ40@ �O�_{F�X_Q\LU�_��V:�t-�Q/B� 1@�Oo!h�&4h+oaG So=oKoyo�o�o?o�o �o�o�o	:�oY@s]k��]4�#&�`�q�%	V3.{00t#mt7H@��*�s$!#�.�� E��qE����E�]\E���HFP=F��{F*HfF@�D�FW�3Fp�?F�MF����F�MF���F�şF���F�=F����G�G�.?�CW�RD�3l)D��E�"��Ex�
E���E�,)F�dRFBFHF�n� F��F���MF�ɽF��,
GlG�g!G)�G�=��GS5�G�iĈ;��
;W�o�|& : E@_z-/�%�#&�)�?�0�&[�B-E�STPARS  �(h L#HR~�A�BLE 1])� G�##i�>� (� �i�i�i�"'T*!i�	i�
i�i�T��#!i�i�i����RDI��g!���ɟ۟����y�O ����������ӯ宙�	S�e# C�����ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��B-~���f"��=�&� 8�J�\���,�>�P��b���#�NUM  ��g!� �+  ��t���_CF�G ���!@�O IMEBF_T�T����e#��N�VE�80t�O�d�N�R {1�� 8 ��#" �� �H�  ����������� '�9�K�]�o������� ��������6#l@GYo}��AN���V;MD���� %7IV_I8]oIINT��bIT��� Bf�8	//�
_TC=/O/�I$��w/�/�RQH�/�/��_�{�@���{�MI_CHA�NZ� �� (3DB/GLVLZ���z��+0ETHERADW ?��~0�)���/�/�?�?s�+0R�OUTx�!
�!��4�?�<SNMA�SKs8��1255.9E�7OIO[O��{�OOLOFS_�DI���%]9OR�QCTRL ���*��MT�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo-l��OPo?otox�PE_�DETAIQ8�JP�GL_CONFI�G �ᄀ�/cell/$�CID$/grp1xo�o $6���?as���� J����'�9�� ]�o���������F�X� ����#�5�G�֏k� }�������şT���� ��1�C�ҟ�y��� ������ӯG�}h�	� �-�?�Q�c���eo��j��g���ҿ���� �a�>�P�b�tφϘ� 'ϼ���������(� ��L�^�p߂ߔߦ�5� ������ ��$��H� Z�l�~����C��� ����� �2���V�h� z�������?������� 
.@��dv� ���M�� *<�`r�������`�Us�er View ��i}}1234567890�/!/�3/E/W/_$� �c/���2�\�/�/�/@�/	??z/�/�3�/ i?{?�?�?�?�?"?�?�.4X?O/OAOSOeOwO�?�O�.5O�O�O��O__+_�OL_�.6 �O�_�_�_�_�_�_>_ o�.7t_9oKo]ooo �o�o�_�o�.8(o�o �o#5G�ohnr� lCamera��o�� �����E�1� C�U��o���������ɏ�I  �v�)�� +�=�O�a�s������ ���ߟ���'�9�`��vW9П������ ��ͯ߯����'�r� K�]�o�������L�^� I<����'�9�K� �oρϓ�޿������ ����߸�^�勪�_� q߃ߕߧ߹�`����� �L�%�7�I�[�m�� &߈usY��������� �#���G�Y�k���� ������������^�'i ��5GYk}�6� ���"�1 CU��^��i��� �����/1/C/ �g/y/�/�/�/�/hz9M/??&?8?J? \?/m?�?�?K/�?�?@�?�?O"O4O�j	�u0�?oO�O�O�O�O�O p?�O�O_�?5_G_Y_ k_}_�_6OHO�p�{3_ �_�_oo0oBo�Ofo xo�o�_�o�o�o�o�o �_�u���oTfx ���Uo���A �,�>�P�b�t�UE h����ҏ����� �>�P�b��������� ��Ο������Իw�,� >�P�b�t���-����� ί����(�:�L� 󟙅@�㯘�����ο �򿙯�(�:υ�^� pςϔϦϸ�_����� O���(�:�L�^�� �ߔߦ��������� �x�$���  �� S�e�w��������������    )�1�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/܋/�  
��( � �G�( 	 �/�/�/�/�/?? =?+?M?O?a?�?�?�?�?�?�*9� � s�$O6OHO��lO~O�O �O�O�O��O�O__ [O8_J_\_n_�_�_�O �_�_�_!_�_o"o4o FoXo�_|o�o�o�_�o �o�o�oeowoT fx�o����� �=�,�>��b�t� ������������� K�(�:�L�^�p���ɏ ۏ��ʟܟ#� ��$� 6�H�Z���~������ Ưد���� �g�D� V�h���������¿Կ �-�?��.�@χ�d� vψϚϬϾ������ �M�*�<�N�`�r߄� �Ϩߺ�������� &�8�J�ߣ߀��� �����������"�i� F�X�j���������� ����/�0w�T�fx������0@� ������� ��#frh�:\tpgl\r�obots\m1�0ia;_7l.xml�_q��������/.��/8/J/\/n/�/�/ �/�/�/�/�/�//? 4?F?X?j?|?�?�?�? �?�?�?�??O0OBO TOfOxO�O�O�O�O�O �O�OO_,_>_P_b_ t_�_�_�_�_�_�_�_ 	_o(o:oLo^opo�o �o�o�o�o�o�oo�o $6HZl~�� ����� �2� D�V�h�z��������ԏ���P ��%<< #?���;���3� U���i���������� ՟�	�7��?�m�S��e��������������$TPGL_OUTPUT � � #�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ������#����2345678901�� ��1�C�U�]����� �ߖߨߺ�����v���@�&�8�J�\���}f� ��������n��� �0�B�T�f���t��� ��������|���, >Pb����� ���� (:L ^p~���� ���$/6/H/Z/l/ ~//�/�/�/�/�/�/ �/
?2?D?V?h?z?? $?�?�?�?�?�?
O�? O@OROdOvO�O O�O��O�O�O�O_�O��} �<_N_`_r_�_�_�]�@��_�_#� ( 	 ��o o6o $oZoHo~olo�o�o�o �o�o�o�o D2 Tzh����� ���
�@�.�d�����2�l�������ҏ 䏾����ʅ�K�]� ��i���m��ɟ۟9� ߟ�����G�Y�3�}� ���w�ů_������ �1�C���+�y���%� ������Ϳ��U�g�-� ?�ٿG�u�O�aϫϽ� ����ύ���)��� _�q���yߧ�Aߓ��� �����%���[�m� ���}����7��� �!���E�W�1�C��� ��������o����� ��AS��W�#u ����e�= �)s�_�� ��/�'/9//E/ o/���/�/Q/�/�/ �/�/#?5?�/Y?k??�W?�?{?�?�?�?{���$TPOFF_L�IM ���@|����ABN_S]V@  �TJ�P_MON �x�D�@�@2��UASTRTCHOK x�F9_�"BVTCOMPA�T/H�AFVWVA/R OM�H3D� �O �O@�bBA_DEFP�ROG %~I�%CL(PSCA�RGA_COVE�YOR_"B_DISPLAY@~N$R�INST_MSK�  v\ `ZI�NUSETP�O$RL�CK�\[QUIC�KMEN�_fTSC�RE�Px��BtpscfT�Q`hiB,`_0iST�J�IRACE_CF�G OI�D�@	�D
?�whHNL 23ZX��a�K 	R�o�o�o�);M_zyeITE�M 2�k ��%$123456�7890��u  �=<����s  #!��{P�?� �C�`��������� �0���T��x�$�J� Џ��ҏ������,� ؟���t�4������� 6�������į(�ЯL� ^�p���B���f�x�ܯ �� ��ۿ6���Z�� ,ϐ�Bϴ�Ϗ�꿪� Ϻ�����V���zό� �����nߔߦ�
��� .�@�R����߈�H�Z� ��f����߽����<� ���r�$����q��� �������H�8�J�\� v�������Pv��� �"4�X* <�H���l� ��T�x�S/ �n/��/�//�/,/ ~/?b/"?�/2?X?j? �/v?�/??�?:?�? OO�?BO�?�?�?NO fO O�O�O6O�OZOlO 5_�OP_�Ot_�_�O�_P_ _�_udS�b�o>�Z�  jr�Z� �aEo<Y
 �Roxo_o�ojUD�1:\�l�� aR_GRP 1�{�� 	 @ EP�o{�o&J8n\~�~p��zhq�o�����u?�   ���>�,�b�P��� t���������Ώ���(��L�:�\���	�U�����SSCB ;2 
k ��� ��*�<�N�`�r�����\UTORIAL� !
k�oϯ�WV�_CONFIG "
m�aBo�o.�ޭ�OUTPUT y#
i���:� ~�������ƿؿ��� � �2�D�V��k�~� �Ϣϴ����������  �2�D�V�g�zߌߞ� ����������
��.� @�R�c�v����� ��������*�<�N� `�q������������ ��&8J\m� �������� "4FXi|� ������// 0/B/T/f/w�/�/�/ �/�/�/�/??,?>? P?b?s/�?�?�?�?�? �?�?OO(O:OLO^O o?�O�O�O�O�O�O�O  __$_6_H_Z_l_� �i��_�_�_�_�_o o(o:oLo^opo�ouO �o�o�o�o�o $ 6HZl~�o�� ����� �2�D� V�h�z������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϟ����� ��������0�B�T� f�xߊߛϮ������� ����,�>�P�b�t� ���߼�������� �(�:�L�^�p�����>wX������� ������_&8J \n������ ���"4FXj |������� /0/B/T/f/x/�/ �/�/�/�/�/�//? ,?>?P?b?t?�?�?�? �?�?�?�??O(O:O LO^OpO�O�O�O�O�O �O�O _O$_6_H_Z_ l_~_�_�_�_�_�_�_ �__ o2oDoVohozo �o�o�o�o�o�o�o	o .@Rdv�� ������*� <�N�`�r��������� ̏ޏ����&�8�J� \�n���������ȟڟ������$TX_�SCREEN 1}$�����}��Q�c�u�������?���>���� �!�3�E���ί{��� ����ÿտL���p�� /�A�S�e�w��� ���������ߐϢ� O�a�s߅ߗߩ� ��� D�����'�9�K��� o��ߓ��������� d�v�#�5�G�Y�k�}� ���������������C�$UAL�RM_MSG ?5-��:� ;� u����� � #)ZM~q�~VSEV  d��TECFG� &-�7� � �@�  A�!   B��
 ��-�7/I/[/ m//�/�/�/�/�/�/��'�GRP 2'�� 0�	 �!/C?V I_BBL�_NOTE (��T���l�2���V2D_EFPRO` %d (%��?��? �?�?O�?,OOPO;O�aO�OqO�O�O�OL<F�KEYDATA �1)-�-0p ��0?3_E__i_{_RZ,(�_�_��POINT 06�_~�_ ANCEL�_�o�PELD_PT�oo!`XT ST�EP:o=oOUCH�UVo�o�QRE INFO�o�o�o�o�o �o,>%bI������� ���/frh/�gui/whit�ehome.pn�g�1�C�U�g�y���  �point������я�����F�RH/FCGTP�/wzcancel��6�H�Z�l�~���arcweld%����ɟ۟���
��nex��;�M�_�q������touchup�+���ѯ�����/info��B�T�f� x���������ʿܿ�  �ϡ�6�H�Z�l�~� ��ϴ���������� ��2�D�V�h�zߌߞ� -���������
��� @�R�d�v���)�� ��������*��/� V�h�z����������� ����
.��Rd v���;��� *<�`r� ���I��// &/8/�J/n/�/�/�/ �/�/W/�/�/?"?4? F?�/j?|?�?�?�?�? S?�?�?OO0OBOTO �?xO�O�O�O�O�OaO �O__,_>_P_�Ob_ �_�_�_�_�_�_o_o@o(o:oLo^o�{kk��������o�o�m�o�o�o�f, ��A(ew^ �������� +��O�6�s���l��� ��͏�����'�� K�]�<���������ɟ ۟�_���#�5�G�Y� k���������ůׯ� x���1�C�U�g��� ��������ӿ����� �-�?�Q�c�u�ϙ� �Ͻ������ς��)� ;�M�_�q߃�ߧ߹� ��������%�7�I� [�m��������� �������3�E�W�i� {�������������� ��/ASew� �r�����  =Oas��� 8���//'/� K/]/o/�/�/�/4/�/ �/�/�/?#?5?�/Y? k?}?�?�?�?B?�?�? �?OO1O�?UOgOyO �O�O�O�OPO�O�O	_ _-_?_�Oc_u_�_�_ �_�_L_�_�_oo)o ;oMo�_qo�o�o�o�o �oZo�o%7I �om�����ڰ �{�� �����(� �J�\�6�,H���@����� Տ�Ώ��/�A�(� e�L������������ ��ܟ� �=�$�a�s� Z���~���ͯ��� �'�9�K�Zo����� ����ɿۿj����#� 5�G�Y��}Ϗϡϳ� ����f�����1�C� U�g��ϋߝ߯����� ��t�	��-�?�Q�c� �߇���������� ���)�;�M�_�q� � ������������~� %7I[m� ������!3 EWi{
��� ���/�//A/S/ e/w/�/��/�/�/�/ �/??�/=?O?a?s? �?�?&?�?�?�?�?O O�?9OKO]OoO�O�O �O4O�O�O�O�O_#_ �OG_Y_k_}_�_�_0_ �_�_�_�_oo1o�_ Uogoyo�o�o�o>o�o �o�o	-�oQc u����L�� ��)�;��_�q��� ������H�ݏ����%�7�I�  K��>  ���t��� ��p���̟��,���� ��!��E�W�>�{�b� ������կ������ /��S�e�L���p��� ��ѿ�ʿ��+�=� /a�sυϗϩϻ�ʏ ������'�9�K��� o߁ߓߥ߷���X��� ���#�5�G���k�}� ��������f���� �1�C�U���y����� ������b���	- ?Qc������ ��p);M _������� �~/%/7/I/[/m/ ��/�/�/�/�/�/z/ ?!?3?E?W?i?{?R� �?�?�?�?�?�? ?O /OAOSOeOwO�OO�O �O�O�O�O_�O+_=_ O_a_s_�__�_�_�_ �_�_oo�_9oKo]o oo�o�o"o�o�o�o�o �o�o5GYk} ��0����� ��C�U�g�y����� ,���ӏ���	��-� ��Q�c�u�������:� ϟ����)���M��_�q����������0�����0��������*�<��,(�m� ϑ�x���ǿ ���ҿ�!��E�,� i�{�bϟφ����ϼ� ������A�S�:�w� ^ߛ߭ߌ?������� �+�:�O�a�s��� ���J�������'� 9���]�o��������� F�������#5G ��k}����T ��1C�g y�����b� 	//-/?/Q/�u/�/ �/�/�/�/^/�/?? )?;?M?_?�/�?�?�? �?�?�?l?OO%O7O IO[O�?O�O�O�O�O �O�O��_!_3_E_W_ i_pO�_�_�_�_�_�_ �_�_o/oAoSoeowo o�o�o�o�o�o�o�o +=Oas� �������'� 9�K�]�o�������� ɏۏ������5�G� Y�k�}������şן ������1�C�U�g� y�����,���ӯ��� 	����?�Q�c�u��� ��(���Ͽ���ϴ)� P+�� P���T�f�x�P��Ϭφ�,���ϐ�� ��%�7��[�B�ߑ� xߵߜ���������� 3�E�,�i�P��t�� ����������OA� S�e�w����������� ����+��Oa s���8��� '�K]o� ���F���/ #/5/�Y/k/}/�/�/ �/B/�/�/�/??1? C?�/g?y?�?�?�?�? P?�?�?	OO-O?O�? cOuO�O�O�O�O�O^O �O__)_;_M_�Oq_ �_�_�_�_�_Z_�_o o%o7oIo[o2�o�o �o�o�o�o�_�o! 3EWi�o��� ���v��/�A� S�e����������я ������+�=�O�a� s��������͟ߟ� ���'�9�K�]�o��� �����ɯۯ����� #�5�G�Y�k�}���� ��ſ׿���Ϝ�1� C�U�g�yϋ�ϯ��� ������	ߘ�-�?�Qߠc�u߇ߙ�p`��}�p`�����@������
����,� M� �q�X������ �������%��I�[� B��f����������� ����!3W>{ �lo����� �/ASew�� *����//� =/O/a/s/�/�/&/�/ �/�/�/??'?�/K? ]?o?�?�?�?4?�?�? �?�?O#O�?GOYOkO }O�O�O�OBO�O�O�O __1_�OU_g_y_�_ �_�_>_�_�_�_	oo -o?o�_couo�o�o�o �oLo�o�o); �o_q����� ����%�7�I�P m��������Ǐُh� ���!�3�E�W��{� ������ß՟d���� �/�A�S�e������� ����ѯ�r���+� =�O�a�𯅿������ Ϳ߿񿀿�'�9�K� ]�o����ϥϷ����� ��|��#�5�G�Y�k� }�ߡ߳��������� ���1�C�U�g�y�� �����������	��p����p���4�F�X�0�z���f�,x��p���� ��;"_qX� |�����% I0mT��� �����!/3/E/ W/i/{/��/�/�/�/ �/�/?�//?A?S?e? w?�??�?�?�?�?�? O�?+O=OOOaOsO�O �O&O�O�O�O�O__ �O9_K_]_o_�_�_"_ �_�_�_�_�_o#o�_ GoYoko}o�o�o0o�o �o�o�o�oCU gy���>�� �	��-��Q�c�u� ������:�Ϗ��� �)�;�/_�q����� ������ݟ���%� 7�I�؟m�������� ǯV�����!�3�E� ԯi�{�������ÿտ d�����/�A�S�� wωϛϭϿ���`��� ��+�=�O�a��υ� �ߩ߻�����n��� '�9�K�]��߁��� ��������|��#�5� G�Y�k���������� ����x�1CUhgyP�{�P�����������,�-� Q8u�n��� ��/�)/;/"/_/ F/�/�/|/�/�/�/�/ ??�/7??[?m?L� �?�?�?�?�?�?��O !O3OEOWOiO{O
O�O �O�O�O�O�O�O_/_ A_S_e_w__�_�_�_ �_�_�_o�_+o=oOo aoso�oo�o�o�o�o �o�o'9K]o ��"����� ��5�G�Y�k�}��� ���ŏ׏����� ��C�U�g�y�����,� ��ӟ���	����?� Q�c�u��������?ϯ ����)�0�M�_� q���������H�ݿ� ��%�7�ƿ[�m�� �ϣϵ�D�������� !�3�E���i�{ߍߟ� ����R�������/� A���e�w����� ��`�����+�=�O� ��s�����������\� ��'9K]�� ������j� #5GY�}�������$U�I_INUSER  ���
!��  ���_MENH�IST 1*
%�  (�  '/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,71,1)/�/�/�/�/� �.c/u%edi�t�"IR_A_HOME�/$?6?H?j�5�/�.CAPTU�RA_CONVEYOR?�?�?�?q�3k?�.DESCA�RGA  DEX,A9�?3OEOWOq)�?u.163�/�O�O�O0�Ovb/�O98�O-_�?_Q_c_f?�?�2L_@�5O�_�_�_l8{_6�_L_FCO�3�_0GoYokot��t^! �a�o�o�o�o�o�o�o �o0BTfx ������� �,�>�P�b�t���� ����Ώ������(� :�L�^�p�������� ʟܟ� ����6�H� Z�l�~���{o��Ưد ���� �#�D�V�h� z�����-�¿Կ��� 
�ϫ�@�R�d�vψ� �Ϭ�;��������� *߹�N�`�r߄ߖߨ� 7���������&�8� ��\�n���� �������"�4�F�I� j�|���������S��� ��0B��Sx �����a� ,>P�t�� ���]�//(/ :/L/^/��/�/�/�/ �/�/��u/?$?6?H? Z?l?o/�?�?�?�?�? �?y?O O2ODOVOhO zO	O�O�O�O�O�O�O �O_._@_R_d_v__ �_�_�_�_�_�_o�_ *o<oNo`oro�oo�o��o�o�o�o�+�$�UI_PANED�ATA 1,����3q � 	�}  f�rh/cgtp/�flexdev.�stm?_wid�th=0&_height=10cp�Tpice=TP&�_lines=1�5&_colum�ns=4cpfon�t=24&_pa�ge=whole�Tp�&)  rim��  Dp�� �(�:�L��^���i� ����ʏ܏Ï ��$� 6��Z�A�~���w�����&� �  }� '�� ���'�9�K���o� �������ɯۯ�T� �#�
�G�.�k�}�d� ����ſ׿������1��U�șs�5s�� �ϧϹ�������B�� ��7�I�[�m�ߑ��� ���߮������!�� E�,�i�P������ ������l�~�/�A�S� e�w������ ����� ��+=��aH �l����� �9 ]oV� ������/#/ vG/Y/��}/�/�/�/ �/�/>/�/�/?1?? U?<?y?�?r?�?�?�? �?�?	O�?-O��p/ uO�O�O�O�O�O"O�O f/_)_;_M___q_�O �_�_�_�_�_�_o�_ %ooIo0omoofo�o �o�o�oLO^O!3 EWi�o� _�� ������A�(� e�L������������ ��܏� �=�O�6�s� �o�o����͟ߟ�� V�'�9��]�o����� �����ۯ¯����� 5��Y�k�R���v����ſ���пπ���}��W�i�{ύϟϱ�)E���I�����&� 8�J�\��π�gߤߋ� ����������"�4�� X�?�|��u��B�������$UI_PO�STYPE  ���� 	� �����QUI�CKMEN  �������RESTORE 1-���  ���K������K�m������+ ��Oas��:� �����"4 �o����Z� ��/#/5/�Y/k/ }/�/�/L�/�/�/D/ ??1?C?U?�/y?�? �?�?�?d?�?�?	OO -O�/�?LO^O�?�O�O �O�O�O�O�O_)_;_ M____�_�_�_�_�_ vO�_�_�_n_7oIo[o moo"o�o�o�o�o�o �o�o!3EWi#�oSCRE3�?8�u1sc��Wu2�t3�t4�tU5�t6�t7�t8�q�sTAT��� xG���USER�pd��rT�p�sks�s�?�4?�5?�6?�7�?�8?���NDO_?CFG .��.��-���PD�q!���None ����_INFOW 1/��ˀE�0%o�B�ԏ��� 9�K�.�o���d����� ɟ۟�������5�����OFFSET 2��ρB�
s}� ����������� ��(�r�,�y�p��� �������ܿ� �J�H�L�:�o�
_ϔ�N��UFRAME  �
t����RTO?L_ABRT��R����ENB����GR�P 13x�D�Cz  A�/�-э� -�?�Q�c�u߇ߙ߫����2�U�ȍ���MS�K  ��ˁ��N6��%É�%�=��%�VCMR�29Nd���p	��� �1: SC�130EF2 *(���
t�I������k�5p��?����@��p���A� 	������x�,��Y�~�T�������A��rm���r B�����q�� e���E�"��F1j U�y�������0��TfO�I�SIONTMOU4�������}y��:SﳸS��� $� FRk:\\��A\k� �� MC�LOG�   oUD1�EX��q' B@ ��2"!,�P/!�T/x/
s � �n6  ���8v/"���`�&�  =����!�
t�  �TRA�IN/�"�"��  �d
3p�)�Z�;d�(�%J=J?X? j?|?�?�?�?�?�?�?@�?OO0OBOw_ �RE�<ل�O�L�EXE�=d���1�-emVMPHA%S�p������P��RTD_FILT�ER 2>d� �L����5_G_Y_k_ }_�_�_�_�_�_G�#_ oo,o>oPoboto�o��o�oM�SHIFT���1?d�
 < ?,+��u�o	B +xOa���� ���,���b�9��	LIVE/S�NAP�vsf�liv�Nt��� ^�U����menu����L��#�����e�@�i	�eMO�A�Nĺ��$W�AITDINEND��؃�O���ߡ����S˟��TIM.������G��� ��;�ʟ������RELE�A�π��<���_ACT��ʨ8���� B�%�xK�����RDIS����ρ�V_AXSR���2C�]�^�V~*1_IR  �F� ��ѿ���� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ���������#�5�G� Y�k�}��������n|XVRf�D�N��$ZABC*21�E�K ,0 2���oZIP�F��O������G�M�PCF_G 1G���04q������H8���S �En@<�P J`u6�Z?�7 �����4�xgyG �= ����������@I]��U�YLI�NDQJ�� ��> ,(  * O/`-EL/�/p/�/�- b�/�/>I/*? �/N?5?G?�?�/�?�? �??�?�?q?&OOJO�1O�?�O�OF�2K��� ����O�L ʳa__:_>�Oj_�>��QA�$SPHERE 2L/-��?�_4O�_�_�_o bOu_Pobo�?�o%oo �o�o�o�o9o(oo �o^�o�i{��o��� ��ZZ� �R�