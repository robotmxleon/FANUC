��   F��A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A #  �����#�AMON_D�O_T   �$PORT_�TYPE  �@NUMJ/SG�NL7 L�$MIN_RAN}GI$MAXr�NOo ALxp V��~ �COUNT>J �AWE08 �� $AWn0ENBJ $�|G1LY_TIV�$WRN_ALM�STP�
�E��C�.�WT�C�
J�AFT_�CHGxAVRG�_INT��{SgAVE�YP1?ER_REG�Tw$WA� SIG�� OP��V/OLTS�����AMP�&AEx �#E_VL� �&D'>% I*f$� _�ANL�  �p 
$US0 S�_CMD � PRIORITY�"�UPPER� $�LOW�$�#$FgDBK�"�RAv ~�!SQ_AVG�#n�#SD_� CE� 8� ��$ �� � �LIN�!$ARC_ENABL�!|� 0DETEC�!~< ELD_SP�$?PD_UNI��!N92DIS�"�ID sIM�#�� � v1WFt2��C�F�" � $�PS_MANUF� �2ODE�L�5PROCES�N0�0WFEEW0EsSC�2�2_FI#1p�1�1�7T _AO�"*�2I�6D�7DC1��6L �"{2 � C�NV� 7   $EQ�zxOD�OU� A<CT�Bd� $?C �2 �?@D�D   , �� MM�!$�D� ��!2 g$F� �BBC�2�NV7	JBSEL�10_NOJDATsA_s@�@ {"�WPpG
{M
�
v�DWP7 L@��L
 �WIR�_CLP4 �L@ASBU8  HG $4���R�4�YPREFx� �U;A_ECU���  JB~ �S �  $BPEtEPf#}!SCH7 � �!��``�1e#dPK*j�FREQ.gULSwbSP�0fg2y��!hyb*g�F�"AI6 �ZCoVG} �hp dD�e�e�`�	�aԤ�dBVB�aZE�ROy}uSLO,]R�`NT�!P�cO	�U\93�L FORM�A0NAra�0J3+	� D�cQWU~XWEIOEX7�4 �A�W�fxccpS_91INp� :1�U�p� �FAUG"t0LO$�0�qP�!�G��R�<�ADp;�STIC|�@�pROBOT��ADY�rERRO&�SE��`S��pƏ!TR��$S�CH�DOG_�@%��0_�ACTIV���I*�C�01�2�q��OTF7 � $
��P��x�nfpNCi0�c ;�f0�*d;�*g0�7f ;�7i0�Fd;�Fg~�Td���TfUP�@�B�sP�CR7�� WGSTK��� =�Hr  ՒƁ%��00��2�X����0A~�3KIPTHE91�S;������PIKEf���0��0WWV�2t�E�_HO;0�0��PH�K-1���� RMT<���SPTL�0p�g$Hz��SW���pd$BBg1_O;NL4�$B�2pf4�bgF�WF�1e2�_R��zE"�!� _W�;6�AND1OFF\���!ND2g�3g��R�S� �A� �SEP�M� | $ �0�@g��e��*f���7b��Ff�TfADA�PT� G�CSEN�S�c��!ݒ��8 � 0?,2���" ��$�1b�!c�7cc� Fa|�Tac�^��'y��&�l��&�!4�&5�&6��"8�W�@�2 HOU��!�o � �SE�0�g4�Q�T<� �6�'��46�q56�0�� %$CURRx7(��"HEATzPe@�!燰"j���i�\p��GAP�#Ti�XPY0��EHP��@��p�DS�@�!GP�0Sf�!$���$GO� 3RI���AM�#/"��#M��jAN3O�BEFB ;�LHV1[5�j��43;1 `H�V�PA�H�r���3��F1��� [@/�SR 7� � 	� RSB �$��0G�m�b�O�J�X��O��DU�IW�"AXQl�2C,1L�"D����?3���8  4�@P֋q]��SGʦ�~�;A8�8 ? $ $�@�CL�$��s	۔��8 $ ;o2� �"��ql��q��� 	PK �P��
��*���q@�Ba��b�@4�5�6:2K�3������FW�q�B<��ALAR���2 ��2�����
�3�Q_R}��
`�.44�F�+�PW,���_@ĸ�Ӕ]� ������Qbwm��t���QDI�c�j��p~pus�R�SIZ���BOAR���1]E7�]�\�h"�0h"��ķ�$V�END��I��DE'VIC��0D�����MAJ��V�#IN`�(�$�uI"�vMA���pFI�0�BW���~�� p $�⠂X�� ⡡��F̀O�R_R��C�^1D4T�O_��O5_R�pR�S<�'�OS�9��U}P� #N� :��0�`�=� �6��6<��9PURG��RKtSTFR�p&���A��.E�.E�AE�D��P-��M%�fMT�����eEM7��Q�5 ���Z$�22�9�P�p���K�p�QADJ�T���NEXT��r_L�E�c��P��X��M ����aA��_�#IV����H�q�2�eFL������P��:����00�8� ��;�WT[𿀻CY��  �aE>�  �	`���`( �bTOTAL!_�Q�c���VI�p�WGWARo��U��A*��PY&1b�uKG@���'" A}�#N�p�  ��SCF�G�1z�LO!O�B:��P�Q�S!x@���GLOB�Pp�⣠� ��NOT�ы$0QI4�*��AVh�Y��$����������e��W_SHFJL�W�X�fkrI�0$�q �e�RY	���p�P��%�ʀLIMS`p�i�@�c7�UIF�e��APCOUPL>�R @ �p�ql��� �qUR�`uN��<�MMYm 0�u0�u�  �����USTOk�    x�0 �qp`� 
@�waEMG�g��1! ,��MGX�Ag���NOzPR ���wa�"� ,/���Ȣ=6Ƞ��3T� )�RT���p�0=����AHER� A�������'"݈{�� �����@���Q�L�� )BD ��2C���7B<�^i3_FIL@�W��7BUG_3SM ���ñF_F����q�, �_4N SV@БTC�P��=Ҕ�DIO��������.a�TM�C��PA�Pq��q�w�x��q�_DYN�V�2Wԣ����KE�YV�GQׂ��F`��?�/B�{�_C��R�TOU���������CAL�Q0�`�� TIp1�P_y�R�T���@��A?2 ��$$CLASS  ������ ��� �-�S�B���  ����IRTUx�����AWAOY1h��[�$�
��K���n�2�f��[�[���g�
�?�������g������� ����(�:�L�^�ppςϑ�l�EXEu� `���������Ͽ�*� <�N�`�r߄ߖߨߺ�\��r@S Rw��� :����#�5�G�Y�k� }���������������l�NLG 2Mx� �����?�ˑ<1�6�`��e��� pp`����{` 2:��)�Ge�neral Pu�rpose��MIG (Vol/ts, 0)���� ����
AWMG�ENL.VR�A*EGLMG19��g�`������ ��'���������������CNV� 2	x��[������ 4aPzUh�� ���//�=/O/ ./s/�/\�/�/b/�/ �/�/?'??K?]?<? �?�?r?�?��E�/�? O�?2ODO#OhOzOYO �O�O�O�O�O�O
__ �?@_R_�Ov_�_g_�_ �_�_�_�_�_o�_(o No�?ro-_�o�o3o�o �o�o�o8J) nM_�{o��� ��� �F�%�j�|� [�������֏�go�� �0�B�!�f�E�W��� {���ҟ������,� >��b�t�������� ί௿�����:�L� +�p����O���ʿU� � �߿$�6��Z�l� KϐϢρ����ϯ��� ߵ�2�D�#�h�z�Y� ��}ߏ��߳���
��NVWP 2|	:i\>�T 
��b��t���USTOM� 2|l  A��������h�	h�d"���DEFSCoH R|�Q��<�b�@Default Schg� ��n��������� ��K"4�Xj �������
)��FBKLOG1 �@��T�῀ � Ugy��12�=O����5L�G_CNT  �����)�IOEX k2�����A ��+C�]$@�������!�
Weld� Spee%��IPM  d$�/�/��/�/??(?:?��O_TF 2��A?��?�?�?�?�?C8=7�����@����?�K)�PCR 2���pI�BH�?��B�C!�FK<D7����>��?�ffAZ �A�"��OFM"@�����/�O@O"@.�����WOELGG��k%*_�F�0�2345678901JRUK%4_y_�_ĝ_HIȩ_7]�OOS�RAM2��IB�$��_oCRGSEL� R<�Q� �	Process# 1oSf2�_ojU3i�o4i�o�5�-mlXS���o7���kn8i'l"@>��� �_);E�s-B� �W�%�Voltage���qsfc%Dw<|!@]y�h����aWire� f�  s�$	 � hc%[&t/�oDS� l*�<�N�`�r����� ����̏ޏ����&��]+zvd"����  ?�#��E�Z"!���a��^/�� ���V���a�aɒCurrent�Amp�=���l �eu���Q�c�u����� ����ϯ����)� ;�M��W���a������ ��	q��)q��Iq��R� ͹ϧg�a�aA��b-� ��-�	q-�)q-�VE!���\e�	q?�����Z�%�������ϻ������PDRuS3 R\zH��jq��C�U�g�����gߩ� ��u߇ߙ������� ��]�o�)�;�M���� �����#������ k�}�7�I�[������� ����1C��I ��Wi���� ��?Q/� �����//)/ ;/M+�U/g){/�/�/�M/�/?cS2�S^=�R��b�S2UPYp�^=�=�o?��33H1>E0=L�S�>I0h!�"��#�$�1t9�g�$q�#?�v�#>�8�8�CWIRE 2�&M<�?�?h�>��3�>�G(=��J*�ESCFG �G�A��Y��OO��E7])COUPL*�0=k
0�vk B`�D�^�L�[�OZW�O��G_�OP_G_Y\�HN�B  ��Ec&FUSTOM  =k�
8ƙy�O&EEMG?OFF !=kS���)BPCR �"�_�@���zqC {sUūMJo�\zt�f_oeo��
Cl�q¨1