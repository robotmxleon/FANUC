��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A   �����
�WVAMP_�T   �$X1  $kX2AY@��/�FC5  �$2ENBA $�DT  / _�R2 d EN�ABLEDnSC�HD_NUMA �SCFG5�� $GROUP��$z ACCEL�@�G$MAX�_FREQ�2 L��DWEL�DE�BUG�PREW�SOUT�P�ULSEASHsIFt 7TYP4�$USE_AE�F} 4$GDO��  f0 �r?�NpWE�AVE_TSK u�V�_GP��SUPPORT_�CFnCNVT_?DONE p }�k}GRP 2�r�� _� �}$� TIME1�to$2'EXT� �(1#&(MODE_�SW�CO3 SW�IT � TPHA|X6  4 � �ECC$�TE�RMNnPEA�Kno!AL O \ � �!I�k$�!N_VSTAR�#!r"���"�%�CYC}L42 
S�� Tv"b $CUR_REL_� ܆!3WPR5 � 
$CEN� �_RI3RADI5U�XIz |] ZIMUTi!�$ELEVAT�IONg5� N�CONTINUOe2xq �MEXAC=�PE�3�6  �H~ �UENCY<A�ITUD4�2�RIGHC�2LE�BL_ANG1 ��OTF_� 	�  $3A�bET��n3C�!$ORGNjHFBKjH��P�q�C��DLDW�H	R�E�_�3�B�C���D�B�C�@�D�A�CCHG�G	Q�F	Q�F	Q�FINC�G=Q�F=Q��F=Q�F�AVCPYC� _T�\#�Y~P#&�@SY��H)@��UPD"0n�$�$CLASS  ����Q��8 <�P�PVERS�1�W�  ����QIRTUAL��_�Q0 2�X��  ��?��@�  HaDae �TWoio{o�o�o`)d�N 2 3k �Hf��uHe@O�Hi�oNc)a� � eG� E`��`9t}
��2  ���=��=�����4s ����jpYq��w�r��Dq��xat ��ujp`��i.�5t8q�q2�b�t����
�9x���� ����̏ҏ���Sb)a�  23k
TDaSI�8� �S����Cph�?m�'����l�D����� Ca��l����k��� ��2�D�V�h�z��l�FIGURE 8��o�v�Hal�f� �������M�(�H� �󈯎�����Ŀֿ�T?CIR1��Pd�}�0�~�h�z�D�Z�l���0�v˜π~����� ��$ߪjN� Hp��4q������@��ʖD�M`g� ���������	��-��?�Q�c�u�`�� �q� �5)�ᐟN`���ᬟ�� ��˟���M�_�q�������������k�Triangle ��z�h߾�M��Ɵ �ύ������/ L� &��g�n��� 	//-/?/Q/c/u/�} DVhz��/�/� �9?K?]?o?�?�?�?�?�?����� O�h ��O2ODOVOhOzO�O �O�O�O�O�O�O
__ .[�?._O"O�_�_�_ �_�_�_�_oo&o8o�Jo\ono�mSCHE�XTENB  �=��ctSTATEw 2�k |o��o�o �gWPR 7�6�L}D�-�_OTF 	8��@)0�q�q���v�)��uAȫs�u@�?  <#�
�?�����mu_GP 2w| ���d�v� ���я㏡+