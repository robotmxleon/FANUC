��  U��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A0  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ���AIO_CNV�w l� RAC��LO�MOD_T�YP@FIR�H�AL�>#IN_O�U�FAC� gINTERCEPf�BI�IZ@!LRM_RECO"w  � ALM�"�ENB���&ONܢ!� MDG/ �0 $DEBUCG1A�"d�$3A�O� ."��!_IF�� P $E/NABL@C#� �P dC#U5K�!M�A�B �"�
� O�G�f d��APCOUPLE, �  $�!PP=_D0CES0�!e8�1�!��R1> Q�� � $SOF�T�T_IDq2TOTAL_EQ� 3$�0�0NO�2U �SPI_INDE�]�5Xq2SCRE�EN_NAM� �e2SIGN�0�e?w;�0PK_FI�0	$THK�Y#GPANE�4 �� DUMMY1"dJD�!UE4RA��RG1R� � _$TIT1d  ��� �Dd�D� �Di@��D5�F6�F7�F8
�F9�G0�G�GPA�E�GhA�E�G1�G �F��G1�G2�B!SB�N_CF�!	 	8� !J� ; 
2L �A_CMNT�?$FLAGS]��CHE"� � EL�LSETUP �
� $HOMEm_ PR<0%�S�MACRO�RREPR�XD0D+�0���R{�T UTOB� U�0 }9DEVIC�CTI�0�� �013�`B�Se#VAL��#ISP_UNI�U`_DODf7{iFR_F�0K%D13���1c�C_WAxqda�jOFF_U0]N�DEL�hLF0pEaA�a7b??a��`$C?��PA#E�C#sATB�d�� oW_PL�0CH/7 <� PU�P��B
2ds�`QgdsD�UT�PHAgpS�F���WELD|H2/0 =Lc�7w7atAING�0�$�r�1�@D2�4%$�AS_LIN;tE��w�t_��2UCC�_AS
BFAIL��DSB"�FAL�0�AB�0�NR�DY��P�z$�YaN�Wq<��`DE6r ��`���+�����tSTK��+�;s7�;sNO�p��[�̈́r��U* Ȁ%�9 � ��  ��q`�G�C�G�+�U�S_FT�vpF�ǂG��SSF��PAUS����ON7xǓHO5U�ŕMI�0�0�ƔSEC�2�ry�i �rHEK0�v8vG#AP�+�	�I� � gGTH���D_I���T= �l���� �`�s9!̅����9!G��UN1���q���#MyO� �cE � �[M�c����RE�V�B7��!XI�� �R  �� OD�P-��dPM� %�;�/�"8�� F�q��
aX�0DfT p{ E RD_E%�~Iq$FSSB�&_$CHKB�pEde#AG� �p�  "
�$Ա� Vt:5���3�Mpa_EDu �� � C2��qS��`�vl �d$OP��0�2�a<�_OK<��Y�TP_C� <�pd�vU �PLAC��^}��p� xaCOM	M� �rD|ƒ��0�`��KO]B BIGA�LLOW� (tK�w�0VAR��xd!�1}!�BL�0S � ,K|a�r�PS�`�0M_O]|=՗�CCG�`=N�! �� ��_I_��� �0�� �B.��1S� ~�CC'BDD�!��I����0�@��84_ CCWp` OOL
��P'�M�M
�n�CHs$MEAdP�d`T�P�!���TRQ�a�CN���FS3��ir�!/0_F��( D�!��v CFfT X0�GRV0��MCqNGFLI���0UJ�p����!� SWIl��&"D�N�P�d��pM~� � �0EED��!��wPo��`�PJedV
�&$�p��1``�P��ELBOF� �=��=�p/0���3P�� ���cẐ�G� �>A0WARNM�`ju���wP��𼠤 CO�R-�8`FLTR^juTRAT Tlp�� $ACC�rT�B� ��r$OR1I�.&��RT�P�p\gMpCHG@I��E3�T{�1�I ̉ra�HK��� �����"�Q���HD(���a�2
BJ{PCT��3�4�5�U6�7�8�9�!����COfS�_rt���3�V�O�LLEC��"MULTI�b
2��A�
1c�O�0T_�R � 4� STY(2�R���).��pp�b�n� |A0@6Kb�Ib$���P�c���UTO=�cE�EXT!Y�
B�!�Q 2 
l��a0��Rpub����  �" ���Q����qc��~#!|��1Y�M�
�P8$  lT}R�� " Lqࠊ/��P��`AX$GJOB׍��W�';IGx# d��? %?78��3�p%���9_MOR��$ et��FN�
CNG&AF�TBA���6䱀JC��9��D@r��1CUR.KPa`/Ek��%��?��ttaoA4��XbJ��_R��|rEC�LJ�r�H�LJ��DA���I�����2G���]QCRfT&�C ��bG����HANC6$LG��iqda��N�*�Ya�Cᇁ�0|rf�R'L±�mTX���nSDB�WnSRA�SnSAZ��P�X��$  ' FCYT��e�_F��Pn�Re�M
P�QIkOh ������1��e����Cg���A���MP�a� ��HK�&AE�Up�p�Q�QI�'�  ]PI���CSXC��Zq( �xs��s��T�R�C�cPN����MG�IsGH"��aWIDR��$VT�P��9�E�F�PA cI�X�P,aQ�1u�CUS�T��U��)R"TI�T����%nAIOV����P_�L����* \q���OR��$!�q���-��OeP��jЅpIp�Q�u��J8�
��0�_�~}pPXWORK��=+�$SK0���nWADBT)PTRw�_ , �l@Ab��s�R0�ؠD��A:0�_C����=�+`H�PL�q��R�A�"��#�D��r�����BJ�b��9�����DB�Q2��-�r~qPR��ΰ�
x ct��. p�E�S�a� �LӉI/��-�( ��0���j� 1%��EsNE���� 2D��b��q	����3H�PC�  .$L��/$Ӄ�����gINE׶�q_D����ROS��E0"2`q��f0�p��PAZ�|tAsbETURN�����MRQ2UA@�C�RŐEWMwp��S�IGN�A&rlPA���W�`0$P�f1$P�P� 	2j���q����!��DQ��f������׶GO_AW;0���pvp��qajDCS'����CYx42O�1P�8�8���2��2��N�@��CtDۣDE�VIѐ 5 P7 $RBֳ���I�P.�i�I_B�Y�q���T�A9�H7NDG�6���x����b�DSBLr3�ͳ��aܢLe7 H �� ���TOFB̶�FE@Бg')��ۣ�f8��cDO�a�� MC9�@�"�`�sr�(��H�P�Wp�X�ܢSLAt4���9IINP!���� ж�ۡ�:D *�SPNp�#�@lƍ�1��W�I1��@J��E�q87�qW�N�NTV#��V n��SKI�STE^�`�b��pڥ�aJ_�Srjb_>���SAF��k���_SVBEX�CLU��po�D�pLX ��YH��%qΉ�I_V9`�bPPLYj���������_ML��L�VR�FY_D��M�IO�`  P�%`�b�Oe��LS�|b��%4}������aP�u���Y�AU NFzf�����)��#"�cD�4Ͱ� S��r�AF� CPX٣e�_� ;j��pTqA#���  ��SGN��<��<@3� P��c_�t�a���qd��rt��`UN>�����<@rD�p]�T`��`��%`����zrEF�p]I>�= @��F��\t6@OTS����|�������孂y Mr�N�IC>2K�GM A���iDAY�sLOCAD���D��5��o�EF pXI�%?j���~cO� �5�_RTRQU�@� D����0Q�p �EԠ��� �?K�%>`� ��GAMP*Pp��A�"�'; DB'��VDUtS�U��CABU�B`�NS9@ID�1WR$�Q!`�V[�V_#� ; ��DI@J$C� �/$VS�SE�#T �BDC�A� ���|�DBf�AE_�;VE�P�0SW!�!�@�x�3�� @�`�O�H�@PP <I	RwqDBB�p�=�!pU����t"BAS�рo'~P�Pn%[�d� B�	� ���RQDWf]%MS� �%AXC'<�;LIFEC���� ��	2N1EB5��D3EBCd@/Ź�Cq`ʡN�4q�6��3OVՐ%6HEh�DB'SUP�1��	2D�_�4j�H1_!C�5š
�7Z�:W�:qa�7�S��"BXZ�PʁEA+Y2HC��T�pސ��NM��zr0P�dgD `L��@HE�VXCSIZ?6k0��[��Nh�UFFI�0���C��������6ܭ�HMSWJEE �8��KEYIMAG�TM���S�A5���F���r��OCVI9E �qF 	�P�LQ�_��?� 	��&`KDG� ��ST��!>R|�FT���FT� FT� FPEMA�ILb �aA|p�FAULSHR�*��;pCOU_��q|pT���U�I< $d�S_�S#�ITճBUFkG�kG@�jpJ`p�0B�Tk�C�p�Rws�PSAV(e �R�+Bd�$ Cg�p��AP/d_ň�$̰_�Pec �iOT�����P@����jA�gAX��sq:p�P��\c_G:3
�YN_e!�pEJ0Df�W�r�d"UMO_0T��F�� �E2���^Јq	K��ey&^�5rH 8)�4��qL���nqL�S�cC_ܐ��K��pu�t��R�A�u�X�nqDSP�FnrPC�{IM5c�s�q�nq��U�w{0�0��PI�PR�nsN!D�@�sT!H��"ûr� Tߑ�s�HSDI�vABSC_�9@`�V��x�v���c~����NV��G ��~�*@�v�PF!�`ad�s0p�a��SC��\��sMER��nqF�BCMP��mpET��⌐M�BFU�0D�U�P?�M�B
�CD�yH��`�S9pR_N)O�ዑN� %�i�Xcg��PSf�C�@%v�C���a~Qd��`U OH����c  d�������}�锍� �9疗疢疮A*�7�8�9�0T��1��1
�1�U1$�11�1>�1K��1X�2f�2���2�
�2�2$�21�2�>�2K�2X�3f�3R�3��
�3�3$�U31�3>�3K�3X�94f��QEXT�TP <sK�p<6p��p2ǋ��QFDR^�QT�PV���b	2p�v�	2REMr�F��0BOVM�sz��A��TROV�ɳDT3`��MX��I�N��Q0�ʶIND����
	�i��`$DG�a{#��4P5�9D���RIV"�=2�0BGEAR�qIO�K��;N0p}ة��(���@�0<Z_MsCM@	1 �F|0;UR"�R ,t� a�? P0�?\��!?��EG ��`a��e�SG � 5P�a�RIM��@��SETUP2_ gT � �STD6� ��<����I�C�`��RwBACrU T[ �RTt)Nz%��+p�IFIQ!+p��А���PT{b[�LU�I1TV � Y�PUR�!�W2�r�<qv��P�� I��$��S��?x#�J�QpCOw`�cVRT|� x$SHO���SASSY��a?5P8�W����A�W�RKFU��15q��25q���*@�X |�N;AV�`��3����*@�R=1��VIS�IJД�SC���EP�c�\�AV��O���B%EX�$PO��I\ ��FMR2b�Y o�X�}p� bpNt�{ߍߟ߶ơP����_f�G�_���B��M4�Y�k�D�GCLFR%DGDMYLD��7�5!6H.�04%�MR�3SZ�@��	 T�FS�`2T[ P!��bs>�`$EX_��B�1�`Ā\2�3�M5��G��9\��
���PWeO�&D�EBUG��"��G�RR�spU�BKUv�O1�� 0PO� ;)' ��' �Mb�LOO�ci!S�M� E7b\$<����� _E ] ��@Y� �TER�M�%^�%[�ORI�Bq� _�%1SM_OpL� `�%^���(�a�&�@UPRbg� -���]�#0^��G:0E�LTO{Q$US]E��NFIc1G2���!���$4_$U;FR��$j�A1�}0=�� OT�7��TqAX�p��3NSTCp�PATM�d@�2PTHJ�;�E4P_bD�H2ARTP`R5�PPa�{RG1REL�:�aS�HFT?�H1�1�8_�N�R�8��& � $�'H@a�q�B���b�SHI@�U�� JaAYLO��a�a����Y�1��~�J�ERVA�3H7�Cp�2�����E����RyC�~�ASYM.q�~�H1WJ[7��E ��1Y�>�U2TCp �a�5�Q=��5P��@���bFORCpMKT�z!:c��'"`&x�0w0�b<�HOb�fd Ԟ2��& X��OCA1E!��$OP����V�t ��#��P��P��`�RŃ�aOUx��3e��R�5Ie h�1���e$PWRL�IM;e�BR_�S�4��� l�3H1UD�_C�R�Bte7�$HSu!^�`ADDR2�H}!AG�2�a�a�a��R��.x�f H!�S��񀌳u��u
�u�S�Ev���!�HS<H�:g $���P�_D�H Y�RrPR�M_��^HTT�P_i�Hx�h (�*�OBJ���b��-$2�LE�3�s��i � #�"�AKB_
�Tp#�rS�P�x���KRL{iHI�TCOUw�B6�L `�rQ��U�`���`SS��JQUERY_FLAQ1��pWR�N1x�jpLgP��PU����O�� �q�!t��/t����<�IOLNw�k�(�� CJq$S�LL$INPU�T_Y$;`��Pt,��C̀SLA� l׀�(�$���C���B1IOgpF�_AShm}�$AL��w��8AِU� �4@_1��݃��情@H�Y1ǧ����a[�UOPen `l�ő2�@�������[`P�c�;`�	������NqU}Ja�o � K�CNEaG4�v7F�Da�֏2J7VpOQR$+J8q�7�I_1z�>��7_LAB�1�Px|���p�APHI���Q{���D�J7�J�-��_KEY�� �K��L�MONx�p�$�XR_���)�WAT�CH_��C��D�E�LD��y����eq� @Р1V�@&�U�C�TR�3U�i��*l��LG��r� -!#�LG�Z�R�`��c��c���FD��I����\!����� �� ��e�Dqf�ce�c�e� ΰe�� e���@0J�_�ѐ1j��qʦ�F �AxǒĞ�Cd(��SB����c��c���ΰ��I�����Ƙ� �ƞ�RS��0 7 (ʀLNe�<sѐ���)��D6Ѽ�UosD��PLM�nC�DAUi�EAwp0���T�u�GH�R1�o�BOOw�t�3 C���`IT\���p� ������SCR��,�㇑DI��Sw0HRGX ���z�d (��o���w�W�o��X�z�JGM^�MN3CHl�n�FN�a��K��PRG��UF���B��FWD��H]L��STP��V�谼 ��Г�RS�HzP��w�CdD��1Rz�: :�^�Unq��9���H�k�����Gw�@( �w�������s�}�OC�/ ��EXv�TUI��I��7�C��O�����<@���	�$��<@��NOA�NAo�A2� VAI̤��tCLUDCS_HI$�!s�1O�
�SI��9S��IGN����ɳ��h�Tc�DEmV<�LL�A�ѧ_BUI �uP��j@T��$��EM@r���]���*"	1vP��j@ހ��~p����1
�2�3�>��� 
0w �C��x�Q@58������IDXa$9 `[����֥1�STƐ�R��Y� <@   /v$E.&C.+�p�mp=&P&����	1x L����`��4@r�`Na�eENwp�dp��?_ y ap7��}p	b���# �MC�7�z �C�CL�DPƐUTRQL�I��TT�94FLAG)"0�Q53�DD��57t�LD55455ORGT�8�H2_ȲF�8�!s�D/r�#�S{ � 	59�455%S�PT0��0y0��4�6RCLMC�D�?�?Iƀ�1pM��p^���|�$D�EBUGGugQDA�TAY��T �U�FE��T)!��M9I6p�T} d@���RQ��0DSTB�`� �F��H�AXR��G�LEXGCES$R>��BMZ`
��~� �B4���BTSq�����F_z@�H�S[�O�H�MwJPTH�� &P�v��r�QMIR� �� � []�R�RCT��N}���VO�ZA�ZL�RC��PC��Q�`D��O��^�CURPX+_THqG�P�`R` |1o)`/d55R^`�`yS�P �B_FR@^�a\fZ_��^ddp�G��* �!KH�� q\��r�Fv$MBu��LI�q�cREQU�IREG�MO�lOX�kfB�$ML� MG�� ap���`|��cZB�ANDU�Sz!�>�5�Z�9sD��Q��IN�p��Q�RSMPf�Sx� �Q�!E]�qRA'qPST� o� 4�LO�Pf�RI ��EX�v�ANG��A�QODkAQG���@$�QG��MFh�������"��%&�2ТfSU�P�%��F `RIG}G�� � ��0 �#1��Ӫ#Q��$$���%#n�א~�א��rPp��wAZw@ETI9��~��Q2�M\p9� �t�pMD�I��) ��� �DA�H�pu���DIA���AN�SW,��w���D���)�!O7��0�Љ+ �QU��VB�70��BL�p�_V@�ъ� �C���sX@�b	|ٰ��P���v����P��KES�!���-�$B����� ND2xFB��2_TX�$�XTRA�1���&�`LO�ЪЋ$RG�&�B�F�8Ҍ|�g��_��rRR2�E��0 #W�e�A�1 d$CALI�@�2�G���2�RI�N����<$R��S�W0"DᣫABC�xD_J��a�����_J3�
�1S�Ps�P��P�-�3P,���?���\�J�hl��2�1O8IM� �2CSKP":��~�$YÛ�J���2Q��̵p��̵·�p_AZ�2�h���ELg�FAO�CMP�s�1!I�R1T�A)�Y�1�i�G�F�1�K�> Y�ZW��SMG�܀�4JG�� SCLP�uSPH_� �0�������=��RTERࠧ��l�IN��ACz�|��� ��r��} _N�я������1hj���?R� �DI��1L�DHP3�����$V��Rs��>$v��p�1�������E�H �$BEL�?w���_ACCEL�0�ث���P_Rـ� ��QT!�*aEX2L6b��3���׀�c��.a�����36cRO
Q_�m�J��P��2�p`��_MG�$DDm�����$FW�0݀�Ӊ�عӤ�~�DE��PP�ABN��RO��EE`���0±�YA(OP��oa_��Y%PaPC��YY���Z�1 �!YN�@A��7����7�M�A��i�g�OL�de�INC a��q����B�����AENCS��Á�B��X���D+`IN"I6bx��ހ��NTVEk�<����23_U���^��LOWL�#0F�0��DF�D�`���� ��`RC����MOS� wT�PP�2��3PERCH  8	OO`�� z�q�! �4!$��!�)b��	A6b�L�tW�����F�
4TRK��!AY[�(cOQI �XM�p/�SQ�� MOMc��BOR�0���D�㣧d��⍠�DU��7bS_BC?KLSH_C�� �@YO`?����*|N�ĵCLALM��p�1�?P6%CHK0|� �GLRTY�� ����Ѕ|1܁_�N'_UMzC�&CzC{ḓ��#��LMT)�_AL�0ú$+��'E�- � �+� ���%��>��C��!4�PC��HI��`q�%C@8�{�.�CN_��N"C�6&��SF�ѯ	V!�p!�����U1��5Y8CAT�.SH����� ?a���X�7aX�L�n�3PA�$��_P�%s_����Pn ��`rD�c%JAaPfC	 OG|s7�TORQU� A�Li���bd����B_W�IU�n��DP_��Ee��EI�KI[Ie�F�P�As�JX��w�VC��0�jS�1q^o��_��wVJRaKq\�R�VDB���M��MPp_DL_��GRV�D�T_��Te��QH_^��S��#jCOS0k1�0hLN�PSktUZd_�Uiv�@Ui'Q�jlEQ�UZN`d�QMY\a�h<b��|Dk�iTHET0$NK23e�rY�]`[CBvCBY�C��ASrqDr'TRq_�Rq�vSB_�pr*uGT	Sֱ��C0��qO�;Cx_Ǧz�c$DU`  ��r����xR�v���1Q��53�NE��7�!I^`q#;��$=�q�Au;�D�"e-h-aLCPH0e����StU ��e���e��f�����f=�V]�VR�O�u�UV��V��V��V��UV��VɋV׉H]�@��|�t��1����H��UH��H��HɋH׉�ON�O]�O�s�O���O��O��O��O*��OɋO�fF�?q�e��P�SPBA�LANCEc�=1LmE�pH_uSP���pf�f�fPFULC������e��{1�+�UTO_[ ��ET1T2_���2NB!�������� �P�p�ҚӞT
O�|���@INSEG�Ҏ=REV��= ��D3IF3�1��1�1�&OB�&!�S°2�@��M!�TLC�HWAR��T�AB�BA�$MECH`Hq�`V�\�q&AXV�P4u�4�@�T�� �
v��Ab���ROB�n CR���j2 ?��MSK_֠��_� P j�_�AR���2����51�2���������$��>�I�Nű�MTCO�M_C\P�Д � h���$N'ORE��Q��.�@�o� 4�@GR�B�a�FLAű$XYZ_DAQ����/DEBU��f�.��mЖ �$/�COD! �҇b���$BUFIwNDX��B_���MOR��� H �����E&��~�^�$޲��o1�� {TA���������G�Ҙ � ?$SIMULp@�����\��OBJE|��\�ADJUSz�m�AY_I�A�D��OUT�@�Ԡ_�_FIb�=��T �@��������q����������D,�FRiI��T�RO�@���E�A�OPW�O�P���,��S�YSBU+���$SCOPT���;!_�U^���PRUN0҅�P�A��D��`�Y� _0��2z��AB��
0^��IMAG!����PϱIM���I�N�P����RGOVCRD�v�e��P����� ��L_R�zA(L�"�0RB� � 1�MC_ED��b� �
0N+�MW	1�MwY191  �sSL����� ����OVSL��SDI5�DEX�3��3
�V�@�N��A��@� ���n�C�0�T��6�_SsET�@��� @�@!��RI^���7_Lq@YLc��\x�0 ���Ta�ޅ@ATUS�$�TRC���ҔB�TM��I��l4p1sU ��� D��!E���4�E�p��� & �EXE�@r!L� "�)�0����UP��!IS��XNN��1l�dQ���PG>՟>L�$SUB���V�ZJMPWAeI�0P��%LO� ���̰[�$RCV?FAIL_C�i��!R��i�r�e1�0�4x���%�`R_PLZ�DBTB�A�2i�B3WD�&Y�UM�@�$�IG�������0TNL�0�$@2R'�T�~@x�@��PPEED5 >�3HADOW�@cÄY�f�E��4�p!D�EFSP�� �# L��|��0_�0���3UNI����0C!IR L�`̰P�%xP1�����Ю@@^Ѻ�� ���X�N�GKETB�@��	@�P42��� h �pSIZE�����ഒ�`ASx�ORZF�ORMATK�*4C�O~ \AǲEMn��|D�3UXC��PsLI%2��� $I�OMP_SWI/�J�E��Wi�Js���P
0%0AL_ !��@�0"�gPBJDpuC�D��$E!��J3D�H� =TV@PDCKC m�>X�CO_J3r�R`QRĢ�	_]���@�C_/1A  � �h�PAY�qҧT�_1�Z2�S�@J3��p�[�U�V�S6�TI�A4�Y5�Y6�MOM�c$cc$cc;�B� ADcHfclHfcPUSpNR)d0uecueb�o �A��ħ` I$PI��Ulq�U*s�Uus �Ujs�UUt�f�kit�t ��v��v_!��m�8��:v3HIG�Cv3 �%�4iv�4�%� ��iv��sxx�!�y�!�%SA�M����tiw�s�%MOV��$�'�
�ް )p%��� #��0�P2� �P%�0�5�`!��@��H��#�INj��@�s q���h��"s�������ӋGAMMǦ���$GET���Є��D�T/�
z�LIB�R9!W2I��$HIB8 _��%�H�E"�bU�AO�r�c�LWJ� ����r���c��Rn�M0��AC50� a ?^I_�p2�/� �B�X�AY��$c/�Hf|��C �$,X� 1���IXR�k�D�>�A!�$@�L�E �8q`���Xq���Z0MSWFL�$M.�@SCRI(7��릀)q�T"@�A����P��UR�$�v��KS_SAVE_�D-B�;#NO�PC `<"�TB�&��_�a�Y W��i�Y�`����pkR#uܸ�SD��p#�s0 �@�,�$�cxY�svY� �x@�<����<!��@}M�ũ � "��YL�c��Y��S ��6�0�� 0����J�@�������	�t�Wq�����`��1�t�M����CL���Q��o� �1T"�@M3�*�� � $��G$WRГ����QR� oTP�vTP�}TP҄T0@���+��C;�@X�0	O~S�AZ�տ@��UԷ� �ՑOMK���V��������̿`C�ON�� / �@�Q_v"� |=Q�B�$i ��c��cB��Z���j�A � CB�����P��P_A��PM� QU�p �� 8@QCOU�M�i�QTH/0HO܋�G�HYS�@ES��F�UE2�8�E@O.�D�  �@P0�@��`UN���q�OVr�а P����%�$��W2ROGRA����2�O����I�T����t�INFOXѱ �A������p�OI� ((�SLEQZv/Nu�/ ����OS��s$�� 4@ENAB|~�� PTIONZ��4(r��4cGCF�l�0J� �A���,�R���CB�OS_ED� �е� �N��K�:�G�E��NUA�UT^�COPY��8 7�1j�MN�NxAE�PRUTfҵ HN� OU�B��0RGADJXѶfTBX_t��2$�0(��мW�P�����v3��#EX� Y�C~��ARGNSrh���ޠLGO���PNYQ_FREQ�bW��MvM!�D��LA��D!�c��@�CRE3�R���IFl�a��NA�q%�$;_G}4TATB0�$>�MAIL�r2��!���B��1�!1�$EL;EMl� �s0vFEASIy@�� �@��2@K�66�V�2�I��0�D"8qJ��L��k2AB�APE��rvpV�!�6BAS&R��52��aU�p��W��$�1�7RMS_TRe3�A���3�ӓp�r�!�4 + !"������	B2 2� ���ԇ�(F�2 'G�2/�_����2SG�gN��DOU��N��!"PRe�m �6G�RID��b�BAR�SZwTYz�"OTIO?`Xѻ���_�$�!��B�DO��i�� � ����PO�R���C�f�BSRV�� )TVDI`�T��P0QCT� MWCpMW4�KY5KY6KY7KY8�/Q�F�l��$VALU�35�(4�w�	�Fh�� !uY����C�!2�F� AN4��R�!R|R!2�TOTAL�s,�a2cPW:#I�AHdREGENFj[b��X�8��R%��V-�T1R�3�rFa_S8��g[`�V���b��2E�#�@L�1�-c7V_H�@DA-��`�pS_Yf���^&S��AR-�2� >�IG_SEC�`dR�%_���dC_�F�Q�E�q�OG6�kjx�SLGEpl�� @>�_%��/�0`9`S���$DE.QU>����s�TE���P�� !�a��aJ�v^�3IL_Mm$;����`��TQ-�6���0Ƨ*��Vh�Cv�P�#1ڀ�M��V1��V1���2��2��3��3
��4��4��$��`ӓ`%�� 0����INA�VIB=�p�]��d�U2`�2l�3`�3l��4`�4l�X�WB�S�B����D $�MC_FP���B%�LC�B�f#cMo�1I��oC ��6���q��KEEP__HNADD�!#�$�0-�C�ѫ C��A⒤�D�O&�"�{���3�D��!a#D�REM[�C�8a�B�������U�$eC�HPWD�  #�SBM�SK�BCOLLAAB/��P@�$a�" �IT$ ��fȕ��� ,(�FL{�W�M�SYNڐ1�M��C`r��G`UP_DLYzX���DELAc��9a�"Y�AD-��z�QSKIPw��� �P��O��NT9�����P_��� ��ҏ�÷�aѹ�ѹ dPкqPк~Pк�PкИPк�Pк9��JS2R ���qX�0TG#r���qr�� �pr����ƐRDCS�W� �_�R�R1�o�=�R�!��J��*D�RGE� T3�ÆBF�LG'����*DSP9C��!UM_r�!�_2TH2NrA<��e� 1� Y���@� 11��� �l����O�v�AT y��.��Q&������@��� *D�Ҙ���H��(�ҥV�2]��c�u�p�ߙ߽߫� U�3]��������(�:� �U�4]�� ]�o����� U�5]���������"��4� U�6]�̀W�i�{�������F�7]��������
.
F�8]��Qcu�ș���S�L�  �1V�p`�L�Z��E%$рpИe)fcIO��Ix�R��POWEC�� M0������U�#d �+��$DSB] � �""c^�QCB��R��M
E�+�R�	D��0E�"���MD"'��M�E� yD�p�'DBG_~@aPD�3%!eaPG
A�@��սS23�2i� ����<P��pICEU�2!`<k$�pARITq!a�OPB�rFLOW>pTR(.b��@�qCU� M%3UX�TA�qINTEORFAC�$��U`����SCHA� t�ݐ"!hpf�$�`�`OM'p�sA���0Iᓴ0Q@IA+ӪTDSv`p���8c3�EFA��p��r�S� k�$�`8b q��R H��6�A ٶ�q  ?2� �S��M ?�	� �$)�s�!0�
eC2`_%pFwDSP)FJOG�`��#�p_P���"ON�g�u���'�	6Ky0_�MIREAb$wpMTY��CAPK�wp4Ц@�4"ASp}@r"At �EBRKH<16=���R�� �B�s�BBP�o0�bC@BSOC�F��NUD1pY1�6��$SVi�D�E_OPGtFSP_D_OVR�k�2�DTRWCORbW� �N�PcVF�@�WB@OVEESF�Z^p�S,r�F�V t'�UFRAv�ZTO�$LCHa��u�2�OVST��B@W Q���BCZ� r&PQ@]s�  @�TIN|�``!$OFSC`C�0@�WD|QdxQ�%Q��E?PTR�!�e"�AFD���AMBS_C��bB5@B<�`�!q�b�a�cSV�� L�k0��s��RG�g�HAMtB_=0�e-b_M�`2�:`OT$CA8@�D�B?pHBKo1~6Tq�IO�cu�pqPPAWz�qhy�t{uu<�:bDVC_W R# �p1��p���Q�u���x-s�u3�v3`��{��0p@SQUR#7@~CAB���,Ӟ`���`��h9�O�`UX~6S�UBCPU�O@S ������dp0ݱ���c��d���$HW_�C]��0ݱrpʆ�8� �Ð�$U��D����ATTRIx�0��O@CYCLw��NECA)��CFLTR_2_FI��/���LP[KC{HKՠ_SCT�CF_�F_�|���FS��b�CHA���d����b�"��RS�DU��Q�3��_�T�hY���c� EM"��M�CT��ݰĀ�����2�DIAG~5RAILAC�sx�M��LO	P7�/V���3� H�3��skPR�pS+� 90қ�C�q&0	,cFU�NC��1RIN����$D����!ʰS	_"@*?p䣸�Mt8���MtCBLȰ����A�
��
�DA`�@�O���LD`0 GPpqw�*A�|�w��TI����AĀ$?CE_RIA��AF��Pn#ò%`ȵ�T2d�C}3�r�aOyI�fDF_LY��Rl1�0LM`#FA>  HRDYO�AM`RG|�Hސ�Q� W�>�MULSE��3���8P�$J_ZJ�zR�W�[FAN_A�LMLV�#��WR=N��HARD�@o6���2$SHADOW `������V����!�Q�E_`s�AU�R��2TO_SBR��6@(�逺s|á@�MPINF8`���S�m�^�REGL���DGy�K�Vm0|��FDAL_N�dsFLۅ9�$Mm��l��g O`L�K�$$Y("V1��2#�� ��CEG[CGP
�A ~/U28S�;���EAXE,GROBn)JRED)FWR  2�A_i�SSY�@D�t�@��S��WRI  �ɀST�*C0�@
nPE�&�w� �""@B��9a��5k�p�OTOn�%`ARY)C�e����[@�FI�@pC$LI�NK�GTH2���0T_��9a%�6�9R[�XYZo2e�7s�OFFA`2� \�LN�uOB'@����0a� h0��FI����0�?T��AD_J �!�2lR?�pq������89R� ��	T�ACL��FDUWb$�9x�TUR��X��z!�bN�X��� )FL[���PH��� |���30�9ROa 1�KN@Ms�/U3��{���8����W3ORQ�6A�����{��@O��N���H�34A��]OV	Ed("M00J��~ ��~��}F1|J�|�{AN��5�~ȱ )!e}@���ve��%��%�6AERSA�	|�E �`��E$A�Ā��ܥ�0�V�S�V�AXc�2 V��ҁ4�%8��)b� �)w��*�*r�*�� �*: �*q �*1� �& ��)��)��)��) ��)��)�9�9��'9D189DEBU��$����0��1Vb�V�ABV�Tq|Q^VIp�� 
B�s�� +E��7G8Q7Gw�7G� 7Gr�7G��7G:7Gq�δF Ȳ4��LAB���)���sGROhB�)��2pB_� ,&��uS��%��FQ*8U�VAND� |�@:$3�_�=!�YW 2q�Z�^�mX�|X5�^�NqT��
c�PVEL����QT��V�SERsVE�P��� $����A�Q!�PPO Hb���`��Q��R�����  $.bTRQK�
 ct�2
`�gȲ2�e��~Q�_ � l����a��ERR��m"Ip� �P�raTOQ���LH�$��f�G�U%H�f���a��	aG� ,�Q#e=`���RA�a 2� �d�b{s�Ta ���$r����"�$ cOCG�p��  dkCOU�NT��` �SF�ZN_CFG	a�# 4ƀ��;�T�Ŀ����3����LsQt��� �(@M��o���`#������uFA���ö�sXd��{�y�aH��S��TO�d�PJ���PHEL��Yr�� 5k�B_B;ASf�RSR�֤�E^�S끐�M�1�g�M�2p�3p�4p�5*p�6p�7p�8�g@��ROO��`9�]�NL��LAB�SN�N��ACKFINpTo���$U��M��� ��_PUV���b�OU�P̠��-��f������&TPFWD_KcARwa��f`RE�T�,�P/�]��QUE����eU �����I ��C-�[�[��Py�[�SEM3A�AAH�An�qSTY�SOސ	�DI�ɠ}s���'���_TM��MANsRQL�[�ENDZ�$KEYSWI�TCH^�s�.�ĔH}EU BEATM��PE�LEvb��@J��Ur�F�s�S3��DO_HOMưOl���EFA PR��Prv����C��O8�<c`�aOV_M����IOCMG˗?�b.�HK��� �DX�׍pU�¹�M�����HFORCΚ�WAR(�)�OM>� � @�4���U��P3�1��2���3��4=� rpOʃ�L����b��UN�LO9����ED���  �SNP�X_ASZr� 0�ЄЍp��$SI=Z��$VAP�e�MULTIP���.�ŰA��� � $H�/����B��S}s�Cr`��FRIFm"pS���������NFO�ODBU ��~P�������UC�N�n��� xU`SI�b�TE�8��SGL*�TA� &opC��C<��+�STMT�\әP��BWe,�S�HOWd�n �SV�7 _G�r� : $�PC�@p7#�!FBZ��P��SPːA�̶��`VD�Оr��� �WaA00 ^T��ɰ��Ӱ��ݰ��T���5��6��7��U8��9��A��B��@���׳A��y���F�ب70���1�1"�1�/�1<�1I�1V�1�c�1p�1}�1��1���1��1��1��2���2�2�2"�2*/�2<�2I�2V�9 T��p�2}�2��2��2��2��2��� `P�>`"�3/�3<�U3I�3V�3c�3p�U3}�3��3��3��U3��3��4k	4�U4�4"�4/�4<�U4I�4V�4c�4p�U4}�4��4��4��U4��4��5k	5�U5�5"�5/�5<�U5I�5V�5c�5p�U5}�5��5��5��U5��5��6k	6�U6�6"�6/�6<�U6I�6V�6c�6p�U6}�6��6��6��U6��6��7k	7�U7�7"�7/�7<�U7I�7V�7c�7p�U7}�7��7��7��7��7��MC��Pz��Ub� `�{@e�
�PV���Q�jU�PR��CM�p��bM�PR9` ��TQ_+pR�P�e(a~��S� `YSL�`�P� � L��jw��A��ؠ; Ѡ�D��VALAUju%�x��A6XF�A�ID_L��^UHI�YZI��$FILE1_L��Ti�$�-���CSAq� h� �pVE_BL�CK���RE��XD_CPU�YM��YA�usȌ_�T�`Y*�F�R �� � PW�-p��<aLAj��SqAcRaKdRUN_FLGde@dhaKd@v�ke�a@d�aKeHF��Wd�`KduATBC2��u� � �B k`(���pĠ���d	�'TDCk`|r�b�p��
u�gTH	�%s�D�1vR��ESERCVE��Rt	�Rt3����`�'p �Xw -$}qLEN��0�t	�}p)�RA���sOLOW_�Ac1}q�vT2�wMO�Q�S���I.��B�Q�y�D�}p�DE���LA3CE,��CCC��B��_MA2��J� ��J�TCVQ�r� �T X�s���������Ѷ�$ ���J+���Mۄ~��Jw������ ��q2��������JK(�VK��:�>��:�sq/�J0O�>�J�JF�JJN�AAL�>�t�F�t�n�4o�5/sX�N1����d�N�
�DL�p_Xќ�*��a�CF6�� `�PG�ROUDPF�Q���N��`C�� �REQUsIR=rؠEBU���yq܆$T�2��6�zp ��$$CL�AF� ���4Z�*�*� O����X�e���~k�IRTUALW��i�AAVM_WR�K 2 ��� 0  G�5a�ͯ٨ʯ.�� ��	��3�*����!�^�E�c���������ɿۿ�㴧�BS�@�� 1�x�� <��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<�~pN�gLMTu�?��7  dQINZl�PPRE_EXEb}� �~AAT��ʖ���IOCNV�Ւ~ �hP�UqS���IO_� w 1��P $����I�4��1��?� ?ܐTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο�����(�:�Q L�ARMRECOV� �c�L�MDG �(BLM_IF m?����� �+���N�`�r߄ߕ�?, 
 �߾߀9�E�������A�NGTOL  ��
 	 A  � Y�k�Q PPLI�CATION ?��� ����ArcTool� �� 
V9.?00P/03j�+�
88340�����F0����161�2�������7D�C3��+��Non}e+�FRA+�� 6�LP_�ACTIV�	�j��UTOMO�D� �Ո	P_CHGAPONL��� ��OUPLE�D 1� � !3��CUR�EQ 1  UT=	==	�������=_�ARC We=l=�AW�ՕAWTOPK�HKY�Dy�9 'EK]o� �����5/�/ #/A/G/Y/k/}/�/�/ �/�/�/1?�/??=? C?U?g?y?�?�?�?�? �?-O�?	OO9O?OQO cOuO�O�O�O�O�O)_ �O__5_;_M___q_ �_�_�_�_�_%o�_o o1o7oIo[omoo�o �o�o�o!�o�o- 3EWi{��� �����)�/�A� S�e�w���������� ����%�+�=�O�a� s����������ߟ� �!�'�9�K�]�o�����OTOC�����DO_CLEAN��|���NM  H���^�p�������A�_DSPDRYRL���HI��<�@M� �&�8�J�\�nπϒ���϶������ψ�MA�X��������
�X��������PLU�GG����
�PRUC˰B:�H�����d�Oi�Կ��SEGF��� ������:� L��&�8�J�\����LAP������ ���������"�4�F��X�j�|�q�TOTA�L,�U�USENU
���� ߨ���O �RGDISPMM�C� ��C���@@M��O���߹RG_STRI�NG 1��
��M��S���
__ITEM1i  n����� ����'9 K]o�������I/O S�IGNALc�Tryout m�odejInp� Simulat{ednOut-,OVERR = 100mIn cycl!%�nProg A�bor7#n$s�tatus�${ c�ess Faul�t�,Aler�$	�Heartbea��#�Hand Broke���/?�?%?7?I?[?m??��e��w�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O__�?WOR��eKQ �?%_s_�_�_�_�_�_ �_�_oo'o9oKo]o�oo�o�o�o�o�nPOc�!�`c[�o$ 6HZl~��� ����� �2�D�8V�h��bDEV�n�� ����̏ޏ���� &�8�J�\�n����������ȟڟ����PALT�=7�c_�_� q���������˯ݯ� ��%�7�I�[�m��8����%�GRI�e ۱O�����'�9�K� ]�oρϓϥϷ����� �����#�5�G�ɿ��R�=��Yߧ߹��� ������%�7�I�[� m�����������m�PREG;�$�� ��K�]�o��������� ��������#5G�Yk}���$A�RG_KPD ?	�������  	]$�	[�]����� SBN_?CONFIG� ��%!$"CII�_SAVE  ��D;� TCE�LLSETUP �
�
%  OM�E_IO��%MOV_H����REP����UT_OBACKs�	�AFRA:\�� ��^'�`� �<(� �M+@ 2�3/04/01 �14:33:48���/�/�/�/-,��?/?A?S?e?w?�?��?�?�?�? �?�?O�?5OGOYOkO }O�O�O,O�O�O�O�O __�OC_U_g_y_�_��_�_�Ё  (!_�#_\ATBCK�CTL.TMP ?DATE.D:��_�oo,o>o#INI�:�o%7#MESSAGS]a^� >hkODE_D�V�7G�eO���o#P�AUS�a!��� ,,		�� ��ow�o- 9;M�q���������;�����d�`TSK  ��m</Bo UPDT̖`[gd���fXW?ZD_ENB[d3��STAZe�����WEPLSCH �R+   b��.�@�R�d�v� ��������П���� �*�<�N�`�r����������̯ޯ����R�ODނ2��4���/��>� % V�{�������ÿտ翀����/�A�SϾWEROBGRP`���r�GWEWEL �2�D���h��� ��'�9�K�]�o߁���ߥ߷��߼	XIS%UN���D��� 	r����@� +�d�O��s���������METER 92b�_ P��&����J���SCRDC�FG 1�N! �[[?� ������������5/�
QW��M_q�� ��2�%�7I���!GR��Р��o��PNAMoE 	��	$n�_EDY`1s��� 
 �%-�PEDT-v��/*/j�� �����.��µ�����/:����%2�/���/a/ ��G(�//?v/�/?�/�#3g?�/�?�/>�?@�?B?T?�?x?�#43O �?�O�?>\O�OO O�ODO�#5�OoOL_�O >(_�_�O�O�__�#6�_;_o__>�__o �_�_No�_�#7�oo �o+o>�o+ro�o��o�#8c/�//� =��>P�t�#!9/��|���=X��Ï
����@��!CR �/�oG�Y�}"���ԏ��|�
���NO_�DEL��GE_�UNUSE��I�GALLOW 1���   (�*SYSTEM�*��	$SERV�_u�.�G�POSREGP�$r�.�G��NUMu�����P�MU���LAY���.�PMP�ALTǧCYC1�0Ԟ�Ѡծ�ULSUǯ���r����L#�\�BOXO{RIy�CUR_I�~��PMCNVæ�I�10����T�4DLIB@�b�	*PROGRAO�PG_MIծ����ALߵ����B<�G�$FLUI_RESU�(u��j������� ������
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� �������������e��LAL_OU�T 6�q#�W?D_ABOR���i�ITR_RTN�  ����l�N�ONSTO���� ��CCG_CONFIG ��7�7���8�����E?_RIA_I����, ���FCFG �����5_LIM^�2�� �� 	n���<j�ߥ�蜀�dPAV�G�P 1?���-?�C��� C�  CU�b�f�b�f��f�b�f0�DZ`�DD���
�����D�v�DZl~�ʆ��x�D/��9�C�M�Wچa��?���HEp��u�"G_P��1� �� d/v/�/�/�/�/�/�HKPAUSf�16�, ���/ ? 6�?L?2?\?�?h?�? �?�?�?�?�?O�?6O�HO.OlO
O9�?��h�COLLECT_9s	`�N�GEN߰��~��B�A�NDE�Cs����1234567890!W��a�pO_1V��
 H+���)l_�_a�k_}_�_ b��_�_o�_�_	obo -o?oQo�ouo�o�o�o �o�o�o:)� M_q�����h��Fm�K �|N�FIO !
Y �A����������ʏb�[TR� 2"F�(��b}�
�؎��#q�x� %[�_MORm$� �)����� ����ǟ���ٛd��*n%r�, %?	!	!I�>���KH���$�R9&�Ow�v�v�C�4  A��
� �x��AA�Cz � B�fPB���Co  @��������:d�
\�I�S'f�\�T_D[EF*� �%�x+�����INUS��&,@�KEY_TOBL  �,v�� �	
��� !"#$%&�'()*+,-.�/*W:;<=>?�@ABC�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~�������������������������������������������������������������������������������͓���������������������������������耇�������������������s��6�d�LCKI�8��d�I�STAs�>��_AUTO_DOr��m���IND�D<�δAR_T1�ϿǃT2�������A�X�C� 2(q�cP8�
SONY X�C-56{�u��U��@���� ���А~�H�R5XY ��߭�R5y7����Aff���6�H� $�m��Z� �����������!����E�W�2�{����T{RL�LETE!���T_SCRE�EN �
�kcsc"UD�MMENU 1)�	?  <u�� 1�:o`CLr �������  &_6H�l~ ����/��I/  /2//V/h/�/�/�/ �/�/�/�/3?
??B? {?R?d?�?�?�?�?�? �?�?/OOOeO<ONO �OrO�O�O�O�O�O_ �O_O_&_8_^_�_n_ �_�_�_�_o�_�_o Ko"o4o�oXojo�o�o �o�o�o�o�o5+���_MANUALH߆�DB9�0�����DBG_ERRL�s*���� >����~uqNUMWLIM����dn��ޠDBPXWOR/K 1+���L��^�p������DBT;B_�� ,�}�����u�RqDB_�AWAY}s͡GwCP n�=����_AL
����yr�YGл�n�nx_�p [1-q�́.��
;�y�z�g�����_MM��IS����@A����ONTIM��M�n��ޖ4�
X��I�MOTNEND�M�H�RECORDw 13�� �����G�O�t�b��� ������į֯m�ޯ� t�)���M�_�q��� ���˿:����%� ��Iϸ�m�ܿ�ϣϵ� ��6���Z��~�3�E� W�i��ύ��ϱ� ��� �����z�/��:��� w�������@��� d��+�=�O���s�^�8l�����Oi�������b�M��sN����8���[���)�;�_JX���W����N/�8�9/�k0.:/q/��/���TOLER7ENC��B�>���L��upCSS_�CNSTCY 2�4,���p�/<�� �/??(?>?L?^?p? �?�?�?�?�?�?�? O�O$O6OHO�$DEV�ICE 25�+ І�O�O�O�O�O �O__+_=_O_���#�HNDGD 6��+ՀCzi^LS 27�Ma_�_�_�_�oo'o9oc_�"PA?RAM 8U�%��duKd�$SLAV�E 9�]nW_C�FG :koKcd�MC:\� L�%04d.CSV�Jo<�c�ofr+"A &sCHp�Q��Kn(*_}g�KfOr|q��zyyq�`JP�Ьsk~<�ρ�lRC_OUT ;�M�ρOo_SGN �<K�4���mE�15-APR-�23 11:32�p�a013�4�:35p�F V�t�g�c�Knd��+�@�S�Þ��j�x�z��cV�ERSION ��V4.0�.1��EFLOG�IC 1=�+ 	�x�`��q���PROG_ENqB)��V2�ULS�� �V�_ACC�LIM����c�q�WRSTJ�Nɐ�3��a�MO�;�uq�b��INIT� >�*K��a OPT�` ?	��Ȓ
 	Rg575Kc�74!�56"�7"�50F�ׄ�L�2"��xp�އ��TO  �z�ů߆]V֐DEX��d&���pݣPATH ;A�A\˯*��<��+HCP_CL?NTID ?�c �{G#|��!�IAG_GRP {2C�i Q�	��ؿÿ��� ���Dϒ�mp1m�10 8901234567n���=�� ?ϜϮω������r������!� 3���\�n����q� Gߩ߻ߙ�����{�� ��9�K�)�o���U� g������������� 3�Y�7�i����+�u� ��������/ gyW��9�� �	�-?�>� �:ϫ����|�@��;/&/_/�˰_O 4Q/�/A/#�/g �/?!?혒$-?W?�/ g?�?o?�?�?m�?E/ O�?ODO/OhOSO�O wO�O�O�O�O�O
_�Op.__R_��<�p c_�_�_C_�_�_ �_�_�_o0o�_@ofo�Qo�ouo�o�o�o��C�T_CONFIG� D��ʓ]��eg�u��ST�BF_TTS��
@J�)s��}�xq<v�p�MAU��?�Q�MS�W_CF�`E�� � ��OCVIE�WPpF�}�a�� ������*�<��� �e�w���������N� �����+�=�̏a� s���������͟\�� ��'�9�K�ڟo��� ������ɯX����� #�5�G�Y��}����� ��ſ׿f�����1�XC�Uϡ|RC�sG]r!�c΍��ϱ������
���.�tSBL�_FAULT �H�ʥxH�GPMS�K2w[��`TDIAOG Iy�qUt���UD1: �67890123C45��x��c�P�o ����*�<�N�`�r� ������������(�;�Vp���@8r��|\��fTRECP����
�ԣ��������� ��1CUgy �������	�0�B�?f�UMP_?OPTION2pT�FaTR�r3sX���PME1uuY_T�EMP  Èϓ3B�Vp��A��UNInp4u����YN_BRK �J��bEDIT�_y�ENT 1K���  ,&�MAIN_SOL?DADURAOP&	G#ON L/P�&IR_HO�ME v/5�&R?EQMENU�/�/�?r��/-?? Q?8?`?�?n?�?�?�? �?�?O�?)O;O"O_O FO�OjO|O�O�O�O�O �O_�O7__[_m_T_��_xY MGDI_�STA��q�%N�C�S1L�{ �P�_�_P
Pd7 Yoko}o�o�o�o�o�o �o�o1CUg y������� �� �.�Fa.�T�f� x���������ҏ��� ��,�>�P�b�t��� ������6������ #�=�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ۟���	��5�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�ӿ����� �-�#�I�[�m��� ������������!� 3�E�W�i�{������� ����������7�A Sew����� ��+=Oa s��������� ///9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?��?�?�?O'/1O COUOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�?�_�_ �_oOo;oMo_oqo �o�o�o�o�o�o�o %7I[m� ��_����o)o 3�E�W�i�{������� ÏՏ�����/�A� S�e�w�������џ ����!�+�=�O�a� s���������ͯ߯� ��'�9�K�]�o��� �����ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߷��� ��������-�?�Q� c�u��������� ����)�;�M�_�q� �����ߝ�������	� ��%7I[m� ������! 3EWi{����� ����///A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?���?�?�?�? /O'O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�? �_�_�_�_Ooo1o CoUogoyo�o�o�o�o �o�o�o	-?Q cu��_���� �_��)�;�M�_�q� ��������ˏݏ�� �%�7�I�[�m��� ����ǟٟ���!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ������� ��'�9�K�]�o�� ���߷���������� #�5�G�Y�k�}��� ������������1� C�U�g�y��ߝ����� ������	-?Q cu������ �);M_q ��y������/ /%/7/I/[/m//�/ �/�/�/�/�/�/?!? 3?E?W?i?���?�? �?y?��?OO/OAO SOeOwO�O�O�O�O�O �O�O__+_=_O_a_ {?�?�_�_�_�_�?�_ oo'o9oKo]ooo�o �o�o�o�o�o�o�o #5GYk�_�� ���_����1� C�U�g�y��������� ӏ���	��-�?�Q� c�}���������ɟ ���)�;�M�_�q� ��������˯ݯ�� �%�7�I�[�u�g��� ����ϟ�����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�m���ߛ߭߿�ٿ ������+�=�O�a� s����������� ��'�9�K���w߁� �������������� #5GYk}�� �����1 CUo�y����� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?gU? �?�?�?��?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_�3_E__? �$EN�ETMODE 1�M�5� W o0o0j5��_�[nPRROR_PROG %{Z�%i6�_�Y�UTAB_LE  {[�?�-o?oQo_g�RSEV�_NUM �R  ��Q�`�Q�_AUTO_EN�B  �U�S�T_;NO�a N{[�Q}�b  *��`���`��`��`�`+��`�o�dHIS�}cm1�P�k_ALMw 1O{[ �j4�li0+�� ����_vb�`  {[�a�R2��nPTCP_VER� !{Z!�_�$�EXTLOG_R�EQ3v�i��SsIZ���STK����e�TOL�  m1Dz;r��A �_BWD��瀠f��R��DI�� P�5���Tm1�STEP�)�;�nPU�OP_D�ȌlQFDR_G�RP 1Q{Y�ad� 	-�ʟ�P����E%�ڭ?��#��[���� �
� ��������!��D� /�h�S���w�������@�ѯ
���.��W
$� ]�fvM�����������B�  �A�  @�33��UO��Ϳ��9�$�F�6 F@]��[�g�"σ�F� ?�  �Ϙ�<P����;O��9 �n���r��������K���/� 舡�[�������[FEATURE R�5���QAr?cTool D�m2�Englis�h Dictio�naryO�4D �Standard�H�Analog �I/OG�AZ�e �Shift��rc� EQ Prog�ram Sele�ct��Softp�ar����Weld���cedures<��@�Core��?�Ramping�۷uto��wa'�U�pdateM�ma�tic Back�upM�{�ground EditE�~R�Camera��=F��Cell�ܠ�nrRndIm�����ommon calib UI��F��sh�����c&��.���neC�.�ty���s����n���M�onitorb�n�tr>�eliab<��N�DHCPD۷��ata Acqu�is���iagn�osw����ocu�ment Vie�we���ua#�h�eck Safesty	�R�han�o Rob��rv��qF
�N�ks" F���(�R�xt we�avx�chJ�xt�. DIO$�nf�iG� endS E�rr��L��s��	r���  �L�F�CTN Menu�; �  TP In�fac(�R�Ge�n��l�Eq L��]��p Mas_k ExcO g��HTJ��xy S�v#�igh-S;peS Ski�����$�mmunic�v�on�Hour�1����Mconun}�2(ncrL�struc�M�KA�REL Cmd.� L�ua�E#R�un-Ti� EnQv;(_�+z�sx��S/WO�Lice�nse5"� Bo�ok(Syste�m)L�MACRO�s,�/Offse�MMR�����MechStop"��t�����%i����6xS ��x�1>od��wit�T8����y.$�r;Optm�?��#��fil"�'g���%ulti-T��E�P�PCM fun4'�9o��6E�^MRegi� r��6ri F
KRF���Nu����nH��Ad�ju�hN�Ҵ٦Mt�atuNA�O
Q�R�DMUot`�scgovei��Eem0�nw��ERZ� ^'ues��9Wo$�_0~N�SNPX b�"vH�SNJCli�}^��urhӝ_z� �%4ujUo� t1ssagE�jU�A�{_bF� U��!n/IK>eMILIB;ob?P Firm^�%n�P1Acc����T�PTX��deln�� XoaA��%&mor�IP Simula(����fu� P]�j���3&��ev.�eV�ri3 �oU�SB po���i�P� a bunexceptS P(Dbu,�uVC�r��8V���rvo�u�[�{�S�PSC�e
�SU�IK�W� �8<�b Pl�FX�Z��� M�#�FQ�uv�n�ԇGrid
Qp�lay΍"`��R2�r.wڊ�RC�g��100iD/14�50��larm �Cause/Pe}dj�Ascii���Load" v�Upl����yc��k"Y@Pp@ %RAp��l��"�NRTL�oS�O�nline Hel���6L�6L@IA��trG�64MB �DRAM��\�FRIOe���tl!�0.L�Gmai#��[�L%�Supmr�1NIР� �cro�LS�U���V�Rmi܉�vrt2SK������W�i� ������̿ÿտ��� �%�/�\�S�eϒω� ���Ͽ��������!� +�X�O�aߎ߅ߗ��� ����������'�T� K�]��������� �������#�P�G�Y� ��}������������� ��LCU�y ������� H?Q~u�� �����//D/ ;/M/z/q/�/�/�/�/ �/�/�/	??@?7?I? v?m??�?�?�?�?�? �?OO<O3OEOrOiO {O�O�O�O�O�O�O_ _8_/_A_n_e_w_�_ �_�_�_�_�_�_o4o +o=ojoaoso�o�o�o �o�o�o�o0'9 f]o����� ���,�#�5�b�Y� k�������Ώŏ׏� ��(��1�^�U�g��� ����ʟ��ӟ���$� �-�Z�Q�c������� Ư��ϯ�� ��)� V�M�_�������¿�� ˿����%�R�I� [ψ�ϑϾϵ����� ����!�N�E�W߄� {ߍߺ߱�������� ��J�A�S��w�� ����������� F�=�O�|�s������� ������B9 Kxo����� ��>5Gt k}�����/ �/:/1/C/p/g/y/ �/�/�/�/�/ ?�/	? 6?-???l?c?u?�?�? �?�?�?�?�?O2O)O ;OhO_OqO�O�O�O�O �O�O�O_._%_7_d_ [_m_�_�_�_�_�_�_ �_�_*o!o3o`oWoio �o�o�o�o�o�o�o�o &/\Se�� ������"�� +�X�O�a��������� ���ߏ���'�T� K�]������������ ۟���#�P�G�Y� ��}��������ׯ� ���L�C�U���y� ������ܿӿ��	� �H�?�Q�~�uχϡ� �����������D� ;�M�z�q߃ߝߧ��� ����
���@�7�I� v�m���������� ����<�3�E�r�i� {������������� 8/Anew� ������4 +=jas��� ����/0/'/9/ f/]/o/�/�/�/�/�/ �/�/�/,?#?5?b?Y? k?�?�?�?�?�?�?�? �?(OO1O^OUOgO�O �O�O�O�O�O�O�O$_�Q  H�541S?Q2DVR�782EW50EUJ�614iW76EUA�WSPQW1�WRC�RuX8�VTU�VJ�545iX�VVCA�MEUCLIO�VR]I�WUIFQV6�W�CMSCh�VST�YLiW2�VCNR�EQV52�VR63�PWSCHEUDOC�VqfCSUEUOR�S�VR869iW0vtW88DVEIOfwR54\VR69�VOESET�W�WJ�Y�WMGEUMASK^EUPRXY5h7EVOC�V�`3�X\V�`�hXgX53�fH^xL�CHvOPLvJ�50HvPS�wMC؋W�p�g55tVMD�SW�w;wOP;wM�PR�Va`0v�`hVP�CMg0��`tW5m0�51�W51P��0�VPRS�g69�0vFRD�VRMC�N)f�hH93hVS�NBAg_wSHL�B)fM߇a`XgNN�lx2hVHTC�VT�MI4fYP�fTPA�fTPTX�EL����p�g8[WYPDVJ�95�VTUT<w9�50vUECvUF]R�VVCC��O�VwVIP4fCSCL�r�`I�xtVWEB�V�HTT�W6WgWImO��CG�IG�oIPGS=�RC4f�HZXR66�VR7��gRN�2HvRjz4�0vu�tV`DVNVD��fD0��F�CTmO�WNN0vOL'h�ENDQVL×SLM�fFVRe XK� ]�o���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ��������� ��1�C�U�g�yߋ� �߯���������	�� -�?�Q�c�u���� ����������)�;� M�_�q����������� ����%7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��� ������)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� =�O�a�sυϗϩϻ����������'� � H541�)�C�2H�R782�I�50I�J614�y�76I�AWSP�Y�1��RCR��8���TU��J545�yܘ�VCAMI�C�LIO�RI�U�IFY�6��CMSyCY��STYLy۽2��CNREY�5�2��R63X�SC�HI�DOCV��C�SUI�ORS��R�869y�0��88�H�EIOh�R54�h�R69��ESE�T�۷�J��WMG�I�MASKI�PRkXY��7I�OC(ꂅ�3��hڅ�x�w�5u3�HLCH��wOPL��J50��PSgMC��u ��{55��MDSW�v��OP��MPR(�p����%�x�PCMH�0����505�1��51X0��P�RSx�69��FR=D�RMCNy���H93x�SNBA�I�SHLBy�MX+���NN(2x�wHTC��TMI���e��TPAh�TPTXi*EL�u �q8g�e�H�J95�ڷTUT��95��U�EC��UFR�V�CC8<O��VIPN��CSC�*��Ii��WEB��HTT���6��WIO�:C�G�;IG�;IPG�S�:RC��Hf�R[66��R7g�RV2��R&4��5@���U�H�NVDx�D0��KF�LCTO��N�N��OLw�END�Y�LG;SLMx�FVRh�(�O_a_s_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �o�o�o�o�o#5 GYk}���� �����1�C�U� g�y���������ӏ� ��	��-�?�Q�c�u� ��������ϟ��� �)�;�M�_�q����� ����˯ݯ���%� 7�I�[�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������ '�9�K�]�o������� ����������#5 GYk}���� ���1CU gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%�}1�STD,�?LANGM�H� `�r߄ߖߨߺ����� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������ 0BTfx��� ����,> Pbt����� ��//(/:/L/^$�RBTL�OPTN�u/�/�/�/�/�+DPNK��/�/??/?M� $�S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_K_]_o_ �_�_�_�_�_�_�_�_ o#o5oGoYoko}o�o �o�o�o�o�o�o 1CUgy��� ����	��-�?� Q�c�u���������Ϗ ����)�;�M�_� q���������˟ݟ� ��%�7�I�[�m�� ������ǯٯ���� !�3�E�W�i�{����� ��ÿտ�����/� A�S�e�wωϛϭϿ� ��������+�=�O� a�s߅ߗߩ߻����� ����'�9�K�]�o� ������������� �#�5�G�Y�k�}��� ������������ 1CUgy��� ����	-? Qcu����� ��//)/;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?m?? �?�?�?�?�?�?�?O !O3OEOWOiO{O�O�O��O�O�O�O�O__�99'U�$FE�AT_ADD ?_	���TQ\P?  	$Xe_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� �����#5�GGTDEMO �RTY    $X������� �///&/8/R/\/�/ �/�/�/�/�/�/�/�/ +?"?4?N?X?�?|?�? �?�?�?�?�?�?'OO 0OJOTO�OxO�O�O�O �O�O�O�O#__,_F_ P_}_t_�_�_�_�_�_ �_�_oo(oBoLoyo po�o�o�o�o�o�o�o $>Hul~ ��������  �:�D�q�h�z����� ��ݏԏ��
��6� @�m�d�v�������ٟ П����2�<�i� `�r�������կ̯ޯ ���.�8�e�\�n� ������ѿȿڿ��� �*�4�a�X�jϗώ� ������������&� 0�]�T�fߓߊߜ��� ���������"�,�Y� P�b��������� ������(�U�L�^� ����������������  $QHZ�~ �������  MDV�z�� �����//I/ @/R//v/�/�/�/�/ �/�/�/??E?<?N? {?r?�?�?�?�?�?�? �?
OOAO8OJOwOnO �O�O�O�O�O�O�O_ _=_4_F_s_j_|_�_ �_�_�_�_�_oo9o 0oBooofoxo�o�o�o �o�o�o�o5,> kbt����� ���1�(�:�g�^� p�������ӏʏ܏��  �-�$�6�c�Z�l��� ����ϟƟ؟���)�  �2�_�V�h������� ˯¯ԯ���%��.� [�R�d�������ǿ�� п���!��*�W�N� `ύτϖ��Ϻ����� ����&�S�J�\߉� �ߒ߿߶�������� �"�O�F�X��|�� ������������ K�B�T���x������� ������G> P}t����� �C:Ly p������	/  //?/6/H/u/l/~/ �/�/�/�/�/?�/? ;?2?D?q?h?z?�?�? �?�?�?O�?
O7O.O @OmOdOvO�O�O�O�O �O�O�O_3_*_<_i_ `_r_�_�_�_�_�_�_ �_o/o&o8oeo\ono �o�o�o�o�o�o�o�o +"4aXj�� ������'�� 0�]�T�f��������� ������#��,�Y� P�b������������ �����(�U�L�^� �����������ܯ� ��$�Q�H�Z���~� �������ؿ���  �M�D�Vσ�zόϦ� ���������
��I� @�R��v߈ߢ߬��� �������E�<�N� {�r���������� ���A�8�J�w�n� �������������� =4Fsj|� �����9 0Bofx��� ����/5/,/>/ k/b/t/�/�/�/�/�/ �/�/?1?(?:?g?^? p?�?�?�?�?�?�?�?  O-O$O6OcOZOlO�O �O�O�O�O�O�O�O)_  _2___V_h_�_�_�_ �_�_�_�_�_%oo.o [oRodo~o�o�o�o�o �o�o�o!*WN `z������ ���&�S�J�\�v� ���������ڏ����"�O�F�r�  i���������П �����*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮��� ��������,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p  qk� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�o, >Pbt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п�����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ���(:L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?h?z?�? �?�?�?�?�?�?
OO .O@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x����� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�\� n��������������� ��"4FXj| �������@0BTfvzm������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o�o�o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n������ ���"�4�F�X�j� |�������ď֏������0�B�T�f�x���$FEAT_DEMOIN  {������~���I�NDEX��������ILECOMP S���ޑ�����ԐSETUP2 Tޕ���  N� �ѓ_AP2B�CK 1Uޙ � �)y�G�V�%=�z�~��h���{� <�ѯ`������+��� O�ޯs������8�Ϳ ߿n�ϒ�'�9�ȿ]� 쿁�ώϷ�F���j� ��ߠ�5���Y�k��� ��߳���T���x�� ���C���g��ߋ�� ,���P��������� ?�Q���u����(��� ��^�����)��M ��q��6�� l�%�2[� ��D�h� /�3/�W/i/��/ /�/@/�/�/v/?�/ /?A?�/e?�/�?�?*? �?N?�?�?�?O�?=O��?JOsO�!�P%�� 2:�*.VRzO�O2@*�O�O/C0�O_E�@PC_H_>2@FR6:3_t^_�_'[T���_�_�]U�_�\���_o FG*.F�OOo1A	_S�=o|lo�o/kST�M�o�o\RbP�o }�o$/kH�oW�gEp�0jGIF����e���-�0jJPG7�a��eM�
�����(ZJS���2@�w�ҏ��%
JavaScript�;�CS�h��fU��� %Casca�ding Sty�le Sheet�s��@
ARGN?AME.DTß&L�`\ן�������ğ�DISP* ���`[���*������H�
TPEINS�.XML˯w�:\�߯����Custo�m Toolba�r �O�PASSW�ORD��$NFR�S:\c�"� %�Password Config�� �?�|��#�YOG�ֿ k�}�ϡ�0�����f� �ϊ�߮���U���y� �r߯�>���b���	� ��-��Q�c��߇�� ��:�L���p������ ;���_������$��� H�����~���7�� ��m��� ��V �z!�E�i {
�.�Rd� �/�/S/�w// �/�/</�/`/�/?�/ +?�/O?�/�/�??�? 8?�?�?n?O�?'O9O �?]O�?�O�O"O�OFO �OjO|O_�O5_�O._ k_�O�__�_�_T_�_ x_oo�_Co�_go�_ o�o,o�oPo�o�o�o �o?Q�ou� �:�^���)� �M��F������6� ˏݏl����%�7�Ə [���� ���D�ٟ h�ҟ���3�W�i� �������ïR��v� �����A�Яe���^� ��*���N������� ��=�O�޿s�ϗ�&� 8���\��π���'߶� K���o߁�ߥ�4��� ��j��ߎ�#����Y��;��$FILE_�DGBCK 1U���F���� < �)�
SUMMARY�.DGc��MD�:�����Di�ag Summa�ry����
CONSLOG�������[���Conso?le log\���	TPACCNQ���%������TP� Account�in}���FR6�:IPKDMP.'ZIP�
'`�����Except�iond��ME?MCHECK��8�����o�Memory Data��;�/YF)	F�TPN�?�C��q�mment T�BDl;�L =��)ETHERNETa������Etherne�t s�figur�a���VDCSV�RF`FXq/��%6  veri?fy allt/>��M+�1%DIF�Fi/O/a/�/� %=�(diff�/�'|�6 CHG01�/��/�/{?�!?�?�"*f992q?X?j?�?
?�?�?@23�?�?�?�O� O�O9FV�TRNDIAG.�LS�O`OrO_���A ��nosti�c_>�T6a)�UPDATES�.MP3_�FRS�:\K_�]��Up�dates Li�st�_�PSRB?WLD.CM�_��wR�_�_p�PS_ROBOWEL�����AHADOW��O�O�O�o�Sh�adow Cha�nges�o=qQbNOTI;/lo�~o�Noti�fic"�o;�+@AG��j�9� ����w���B� �f�x����+���ҏ a��������'�P�ߏ t������9�Ο]�� ���(���L�^�ퟂ� ���5���ܯk� ��� $�6�ůZ��~���� ��C�ؿ�y�ϝ�2� ��?�h�����ϰ��� Q���u�
�߫�@��� d�v�ߚ�)߾�M��� �߃���<�N���r� ���7���[���� ��&���J���W���� ��3�����i�����" 4��X��|�� A�e��0� Tf����O �s//�>/�b/ �o/�/'/�/K/�/�/ �/?�/:?L?�/p?�/ �?�?5?�?Y?�?}?�? $O�?HO�?lO~OO�O 1O�O�OgO�O�O _2_ �OV_�Oz_	_�_�_?_ �_c_�_
o�_.o�_Ro do�_�oo�o�oMo�o qo�o<�o`�o ��%�I�� ��8�J��n���� !���ȏW��{��"� ��F�Տj�|����/� ğ֟e��������+� T��x������=�ү a������,���P�b� 񯆿���9����o� ϓ�(�:�ɿ^��� ��#ϸ�G�����}�����6���C�l�N��$�FILE_FRS�PRT  ���V�������MDONLY� 1U��N� �
 �)MD:�_VDAEXTP.ZZZs�$���
��6%NO �Back fil�e ��N�S�6 �\��߀�Iߍ���� ��i������4���X� j���������S��� w���B��f�� ��+�O��� �>P�t� '��]��/(/ �L/�p/�//�/5/��/�/��VISBC�K�؝���*.V�D�/'?� FR:�\� ION\DA�TA\?�"� �Vision VD(�S?a/�?�?�/�? �/�?�?O+O�?OO�? sO�OO�O8O�O\OnO _�O'_9_�O]_�O�_ _�_�_F_�_j_�_o �_5o�_Yo�_�_�oo �o�o�o�oxo�o C�og�o��,��P�t��{�LU�I_CONFIG7 V��	1&�� $ ���{ ��}�������ŏ׏�e�|x��!�3�E� W�g�����������ҟ i����,�>�P�� t���������ίe�� ��(�:�L��p��� ������ʿa�� �� $�6�H�߿l�~ϐϢ� ����]������ �2� D���h�zߌߞ߰��� Y�����
��.���?� d�v����C����� ����*���N�`�r� ������?������� &��J\n�� �;����" �FXj|��7 ����//�B/ T/f/x/�/!/�/�/�/ �/�/?�/,?>?P?b? t?�??�?�?�?�?�? O�?(O:OLO^OpO�O O�O�O�O�O�O _�O $_6_H_Z_l_~__�_ �_�_�_�_�_�_ o2o DoVohozoo�o�o�o �o�o}o�o.@R d�o������ y��*�<�N�`�� ��������̏ޏu�� �&�8�J�\�󏀟�� ����ȟڟq����"� 4�F�X��|��������į֯f��|�$�FLUI_DAT�A W���>�j����RESULT 2�X�0� ��T�/wiza�rd/guide�d/steps/?Expert�g� y���������ӿ����	��)��Con�tinue wi�th GD�ance)�d�vψϚϬϾ����������*� ��-��I�0� �r�I�	��i��;�ps,ߴ����� ����� �2�D�V�h� z�9�r���������� ����1�C�U�g�y����i�[�m����torch��% 7I[m��� �����!3E Wi{���������������wproc��U/g/y/�/�/ �/�/�/�/�/	??� ??Q?c?u?�?�?�?�? �?�?�?OO)O���DO/����M�Ti�meUS/DST 3O�O�O�O�O__'_�9_K_]_o_2�DisablRϤ_�_�_ �_�_�_o"o4oFoXoTjo|n�j�eO`WOiO{O�O�B24�O /ASew� ���~_�_��� +�=�O�a�s������� ��͏�o�o�o�o��:�~L�RegionЏ _�q���������˟ݟ����.�AmericaI/M�_�q� ��������˯ݯ���.�ہyE���]��1��BEdi��$��� ſ׿�����1�C��U�g�*; Touc�h Panel ��� (recommen��)uϺ��� ������&�8�J�\�n�-��=�O���s���>�Bacces<�� �*�<�N�`�r�������)<Conn�ect to N?etwork�� � �$�6�H�Z�l�~���������1��鏣�����!�ߝ@Int?roductK�^ p�������  -?6HZl~ �������/ / =O��=/�b 0�/�/�/�/�/�/�/ ?#?5?G?Y?k?*�? �?�?�?�?�?�?OO 1OCOUOgO׈@ ]/>G*���~�O�O }/�O�O__*_<_N_ `_r_�_�_�_�_y?�_ �_oo&o8oJo\ono �o�o�o�ouO�O�O�O �O4FXj|� ��������_ 0�B�T�f�x������� ��ҏ������o�o �o_�!��������Ο �����(�:�L�^� ���������ʯܯ�  ��$�6�H�Z�l�+� =�O���s�ؿ����  �2�D�V�h�zόϞ� ��o�������
��.� @�R�d�v߈ߚ߬߾� }��ߡ��ſ*�<�N� `�r��������� ����%�8�J�\�n� ���������������� ��1��U�|� ������ 0BTf%���� ����//,/>/ P/b/!�/E�/ik/ �/�/??(?:?L?^? p?�?�?�?�?w�?�?  OO$O6OHOZOlO~O �O�O�Os/�O�/�O_ �?2_D_V_h_z_�_�_ �_�_�_�_�_
o�?.o @oRodovo�o�o�o�o �o�o�o�O_�O3 ]_������ ���&�8�J�\�o ��������ȏڏ��� �"�4�F�X�a; ����q֟����� 0�B�T�f�x������� m�ү�����,�>� P�b�t�������i�{� �����ß(�:�L�^� pςϔϦϸ�������  ߿�$�6�H�Z�l�~� �ߢߴ���������� Ϳ߿�S��z��� ����������
��.� @�R��v��������� ������*<N `�1�C�g��� �&8J\n ���c����� /"/4/F/X/j/|/�/ �/�/q�/��/�? 0?B?T?f?x?�?�?�? �?�?�?�?O?,O>O PObOtO�O�O�O�O�O �O�O_�/%_�/I_? p_�_�_�_�_�_�_�_  oo$o6oHoZoO~o �o�o�o�o�o�o�o  2DV_w9_� ]__���
��.� @�R�d�v�������ko Џ����*�<�N� `�r�������gɟ� ���Ï&�8�J�\�n� ��������ȯگ��� ��"�4�F�X�j�|��� ����Ŀֿ������ ݟ'�Q��xϊϜϮ� ����������,�>� P��t߆ߘߪ߼��� ������(�:�L�� U�/�y��e�������  ��$�6�H�Z�l�~� ����a���������  2DVhz�� ]�o������. @Rdv���� �����/*/</N/ `/r/�/�/�/�/�/�/ �/?���G?	n? �?�?�?�?�?�?�?�? O"O4OFO/jO|O�O �O�O�O�O�O�O__ 0_B_T_?%?7?�_[? �_�_�_�_oo,o>o Poboto�o�oWO�o�o �o�o(:L^ p���e_��_� �_�$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ������ =��d�v��������� Я�����*�<�N� �r���������̿޿ ���&�8�J�	�k� -���Q�S��������� �"�4�F�X�j�|ߎ� ��_����������� 0�B�T�f�x���[� ���������,�>� P�b�t����������� ������(:L^ p������� ������E�l~ �������/  /2/D/h/z/�/�/ �/�/�/�/�/
??.? @?�I#m?�?Y�? �?�?�?OO*O<ONO `OrO�O�OU/�O�O�O �O__&_8_J_\_n_ �_�_Q?c?u?�?�_�? o"o4oFoXojo|o�o �o�o�o�o�o�O 0BTfx��� �����_�_�_;� �_b�t���������Ώ �����(�:��o^� p���������ʟܟ�  ��$�6�H���+� ��O���Ưد����  �2�D�V�h�z���K� ��¿Կ���
��.� @�R�d�vψϚ�Y��� }��ϡ���*�<�N� `�r߄ߖߨߺ����� ����&�8�J�\�n� ������������ ���1���X�j�|��� ������������ 0B�fx��� ����,> ��_!��E�G�� ��//(/:/L/^/ p/�/�/S�/�/�/�/  ??$?6?H?Z?l?~? �?O�?s�?�?�/O  O2ODOVOhOzO�O�O �O�O�O�O�/
__._ @_R_d_v_�_�_�_�_ �_�_�?�?�?o9o�? `oro�o�o�o�o�o�o �o&8�O\n �������� �"�4��_=ooa��� Mo��ď֏����� 0�B�T�f�x���I�� ��ҟ�����,�>� P�b�t���E�W�i�{� ݯ����(�:�L�^� p���������ʿܿ��  ��$�6�H�Z�l�~� �Ϣϴ������ϩ��� ͯ/��V�h�zߌߞ� ����������
��.� �R�d�v����� ��������*�<��� �߁�Cߨ������� ��&8J\n �?������ "4FXj|� M��q�����// 0/B/T/f/x/�/�/�/ �/�/�/�??,?>? P?b?t?�?�?�?�?�? �?�O�%O�LO^O pO�O�O�O�O�O�O�O  __$_6_�/Z_l_~_ �_�_�_�_�_�_�_o  o2o�?SoOwo9O;o �o�o�o�o�o
. @Rdv�G_�� �����*�<�N� `�r���Co��goɏۏ ���&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��� ����į֯��ߏ��� -��T�f�x������� ��ҿ�����,�� P�b�tφϘϪϼ��� ������(��1�� U��A��߸�������  ��$�6�H�Z�l�~� =Ϣ�����������  �2�D�V�h�z�9�K� ]�o�������
. @Rdv���� ����*<N `r������ ������#/��J/\/n/ �/�/�/�/�/�/�/�/ ?"?�F?X?j?|?�? �?�?�?�?�?�?OO 0O�//uO7/�O�O �O�O�O�O__,_>_ P_b_t_3?�_�_�_�_ �_�_oo(o:oLo^o po�oAO�oeO�o�O�o  $6HZl~ ������o��  �2�D�V�h�z����� ��ԏ�o���o��o @�R�d�v��������� П�����*��N� `�r���������̯ޯ ���&��G�	�k� -�/�����ȿڿ��� �"�4�F�X�j�|�;� �ϲ����������� 0�B�T�f�x�7���[� ���ߓ�����,�>� P�b�t������� ������(�:�L�^� p��������������� ����!��HZl~ �������  ��DVhz�� �����
//�� %��I/s/5�/�/�/ �/�/�/??*?<?N? `?r?1�?�?�?�?�? �?OO&O8OJO\OnO -/?/Q/c/�O�/�O�O _"_4_F_X_j_|_�_ �_�_�_�?�_�_oo 0oBoTofoxo�o�o�o �o�o�O�O�O�O> Pbt����� �����_:�L�^� p���������ʏ܏�  ��$��o�oi�+ ������Ɵ؟����  �2�D�V�h�'�y��� ��¯ԯ���
��.� @�R�d�v�5���Y��� }������*�<�N� `�rτϖϨϺ���ݿ ����&�8�J�\�n� �ߒߤ߶��߇��߫� �Ͽ4�F�X�j�|�� ������������� ��B�T�f�x������� ����������; ��_!�#���� ��(:L^ p/�������  //$/6/H/Z/l/+ �/O�/�/��/�/?  ?2?D?V?h?z?�?�? �?�?��?�?
OO.O @OROdOvO�O�O�O�O }/�/�/�O_�/<_N_ `_r_�_�_�_�_�_�_ �_oo�?8oJo\ono �o�o�o�o�o�o�o�o �O_�O=g)_� �������� 0�B�T�f�%o������ ��ҏ�����,�>� P�b�!3EW��{ �����(�:�L�^� p���������w�ܯ�  ��$�6�H�Z�l�~� ������ƿ������� ͟2�D�V�h�zόϞ� ����������
�ɯ.� @�R�d�v߈ߚ߬߾� ��������׿��� ]�τ�������� ����&�8�J�\�� m��������������� "4FXj)� M�q���� 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/{ �/�?�(?:?L?^? p?�?�?�?�?�?�?�?  OO�6OHOZOlO~O �O�O�O�O�O�O�O_ �//_�/S_?_�_�_ �_�_�_�_�_
oo.o @oRodo#O�o�o�o�o �o�o�o*<N `_�C_��{o� ���&�8�J�\�n� ��������uoڏ��� �"�4�F�X�j�|��� ����q��ߟ	�� 0�B�T�f�x������� ��ү����Ǐ,�>� P�b�t���������ο ���ß��1�[� ��ϔϦϸ�������  ��$�6�H�Z��~� �ߢߴ����������  �2�D�V��'�9�K� ��o�������
��.� @�R�d�v�������k� ������*<N `r����y�� �����&8J\n �������� ��"/4/F/X/j/|/�/ �/�/�/�/�/�/?� ��Q?x?�?�?�? �?�?�?�?OO,O>O PO/aO�O�O�O�O�O �O�O__(_:_L_^_ ?_A?�_e?�_�_�_  oo$o6oHoZolo~o �o�o�o�_�o�o�o  2DVhz�� �o_��_��_�.� @�R�d�v��������� Џ����o*�<�N� `�r���������̟ޟ ���#��G�	�� ��������ȯگ��� �"�4�F�X��|��� ����Ŀֿ����� 0�B�T��u�7��ϫ� o���������,�>� P�b�t߆ߘߪ�i��� ������(�:�L�^� p����eϯω��� ���$�6�H�Z�l�~� ����������������  2DVhz�� ���������� %O�v���� ���//*/</N/ r/�/�/�/�/�/�/ �/??&?8?J?	 -?�?c�?�?�?�? O"O4OFOXOjO|O�O �O_/�O�O�O�O__ 0_B_T_f_x_�_�_�_ m??�?�_�?o,o>o Poboto�o�o�o�o�o �o�o�O(:L^ p�������  ��_�_�_E�ol�~� ������Ə؏����  �2�D�U�z����� ��ԟ���
��.� @�R��s�5���Y��� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ�c��χ��ϫ� �"�4�F�X�j�|ߎ� �߲��������߹�� 0�B�T�f�x���� ������������;� ����t����������� ����(:L� p�������  $6H�i+� ��c����/  /2/D/V/h/z/�/�/ ]�/�/�/�/
??.? @?R?d?v?�?�?Y� }�?�?�O*O<ONO `OrO�O�O�O�O�O�O �O�/_&_8_J_\_n_ �_�_�_�_�_�_�_�? �?�?oCoOjo|o�o �o�o�o�o�o�o 0B_fx��� ������,�>� �_o!o3o��Wo��Ώ �����(�:�L�^� p�����S��ʟܟ�  ��$�6�H�Z�l�~� ����a�s���篩��  �2�D�V�h�z����� ��¿Կ濥�
��.� @�R�d�vψϚϬϾ� �����ϳ�ůׯ9��� `�r߄ߖߨߺ����� ����&�8���I�n� ������������� �"�4�F��g�)ߋ� M߲��������� 0BTfx���� ����,> Pbt��W��{� ���//(/:/L/^/ p/�/�/�/�/�/�/�/ �?$?6?H?Z?l?~? �?�?�?�?�?�?�O �/O��?hOzO�O�O �O�O�O�O�O
__._ @_�/d_v_�_�_�_�_ �_�_�_oo*o<o�? ]oO�o�oW_�o�o�o �o&8J\n ��Q_����� �"�4�F�X�j�|��� Mo�oqo��叧o�� 0�B�T�f�x������� ��ҟ䟣��,�>� P�b�t���������ί ௟��Ï�7���^� p���������ʿܿ�  ��$�6���Z�l�~� �Ϣϴ����������  �2����'���K� ����������
��.� @�R�d�v��GϬ�� ��������*�<�N� `�r�����U�g�y��� ��&8J\n ��������� "4FXj|� ����������� -/��T/f/x/�/�/�/ �/�/�/�/??,?� =?b?t?�?�?�?�?�? �?�?OO(O:O�[O /OA/�O�O�O�O�O  __$_6_H_Z_l_~_ �_�O�_�_�_�_�_o  o2oDoVohozo�oKO �ooO�o�O�o
. @Rdv���� ���_��*�<�N� `�r���������̏ޏ �o���o#��o�\�n� ��������ȟڟ��� �"�4��X�j�|��� ����į֯����� 0��Q��u���K��� ��ҿ�����,�>� P�b�tφ�E��ϼ��� ������(�:�L�^� p߂�A���e����ߛ�  ��$�6�H�Z�l�~� ������������  �2�D�V�h�z����� ���������߷�+ ��Rdv���� ���*��N `r������ �//&/����	 }/?�/�/�/�/�/�/ ?"?4?F?X?j?|?; �?�?�?�?�?�?OO 0OBOTOfOxO�OI/[/ m/�O�/�O__,_>_ P_b_t_�_�_�_�_�_ �?�_oo(o:oLo^o po�o�o�o�o�o�o�O �O�O!�OHZl~ ��������  ��_1�V�h�z����� ��ԏ���
��.� �oO�s�5������ П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��?���c�ſ����� �"�4�F�X�j�|ώ� �ϲ����ϕ����� 0�B�T�f�xߊߜ߮� ���ߑ��ߵ��ٿ�� P�b�t������� ������(���L�^� p���������������  $��E�i{ ?�������  2DVhz9�� �����
//./ @/R/d/v/5Y�/ �/��/??*?<?N? `?r?�?�?�?�?�?� �?OO&O8OJO\OnO �O�O�O�O�O�/�/�/��O_%Q�$FMR�2_GRP 1Y�%U� ��C4  B�.�0	 �0c_u\�`PF�6 F@ �S�Q�T�J`S�_�]`P�?�  �_�_<P��a;O��9' n�e�]A`+o6=kBH]SB�YPX`�;a@�33ce�\x�_�o�Y@UO߯a �o�_�o�o�o�o4 XC|g�����}9R_CFG =ZF[T ���(�:��{NO ^FZ
F0p� u���|RM_CHKTYP  6Q�0NP�PPP8QROM��_�MIN���3��꽀�|`X9PSSB��s[%U aV��5�
����uTP_DEF__OW  �4NS>1�IRCOM��B���$GENOVR/D_DO���1o��THR�� d��d�u�_ENBa� ^u�RAVC?S\Ӈހ ��U"����1��?�P�sj [�ՑOUBPbF\�x�sXF�sU<�� �]ǯq���X���3C�YP�YPa�%��d��1A@M��?�U�vY��#�֐SMT?Sc�RP��4��$HOSTC�rs1dFY߀��?�_P MC�4L��
��6  27�.0Z�1C�  e:χϙϫϽ���uπ�� ��$�G�����	�anonymou�sK�yߋߝ߯��� 	�^P����8�:�'� n�K�]�o����Ϸ� ��������X�5�G� Y�k�}���������� �0���1CU�� y�������,� 	-?Q������ ������// )/pM/_/q/�/�/� ��/�/�/??%?l ~�m?�/�?��?�? �?�?2/O!O3OEOWO z?�?�/�O�O�O�O�O .?@?R?d?fOS_�?w_ �_�_�_�_O�_�_o o+oN_�O�Oso�o�o �o�o__&_:o' n_K]o�Ho>� ����Xo5�G� Y�k�}��o�o�o�o� Ώ0��1�C�U�� y�����������,��	��-�?�Q����E�NT 1e�� sP!ڟ��  ����ï��篪��ί /��;��d���L��� p�ѿ�������ܿ� O��s�6ϗ�Zϻ�~� ���ϴ����9���]�  �Vߓ߂߷�z��ߞ� �������4�Y��}� @��d������������C��g�*�QUICC0t�P�b�����1���������2��c!ROUTERd@R��!PCJOG���!192�.168.0.1�0����CAMPRYT�!�1� +RT}/A��h�NAME !~u�!ROBO��S_CFG 1�du� ��Auto-st�arted��FTP��;!͏ϟf/ ��/�/�/�/�/o��/ ??,?O/=?�/t?�? �?�?�?��/&/8/O L?n/,O]OoO�O�OZ? �O�O�O�O�O"O�O5_ G_Y_k_}_�_������ ʏ_�_BOo1oCoUo go._�o�o�o�o�o�_ xo	-?Qc�_ �_�_��o�o�� �)��oM�_�q����� �:���ݏ���%� l~��������� ǟٟ���ď!�3�E� W�i��������ïկ ���@�R�d�A�x�e� ������������|��� ��+�N�O��sυ� �ϩϻ���&�8�:� �n�K�]�o߁ߓ�Z� ����������"ߤ�5� G�Y�k�}�������� �����B��1�C�U� g�.������������ x�	-?Q��_ERR f��aqPDUSIZW  ��^����>�WRD ?�%���  guest�����);�S�CD_GROUP� 3g, !��� �LOA���RES�T�M� $�T_�ENBs TTP�_AUTH 1h�� <!iPendanGR.����A!KAR�EL:*R/[/m-�KC�/�/�/z V�ISION SE!Tk?�/F!?? 1?w#U?C?m?g?�?�?��?�?�?�>!$CTR/L i�;H���
��FFF9�E3�?��FRS�:DEFAULT�`LFANUC� Web Server`JNB!$�� 	L�O�O�O__,_o�WR_CONFI�G jp�`OqIDL_�CPU_PC@���B����P BH��UMIN�\x�UGNR_IOz������PNPT_SI�M_DO�V�[S�TAL_SCRN��V �6F�QTPM?ODNTOLg�[�ARTY�X�Q�V� �%  gx�SOL_NK 1k�} �o�o�o�o�o �b_MASTE�Pzi��UOSLAVE �l�AuRAMCOACHE0(bO'!O_CFGr�c�s�UO0��rCYC�Lq�uy@_ASG� 1maW�
  �)�;�M�_�q��� ������ˏݏ��{��rNUM��	
�rIPo�wRTRY_CN@�R�
�r�a_UPD��a�b� �r�p�rnP~�u��u�PSDT_�ISOLC  �P{v"�J23_�DSrd.N�OGvg1oP{<��sd<�P� ?��DR��?��館Q�� ̯ޯ𯯯�&�8�J�������*��P�qi���PhpECso�UK_ANJI_*pK�_�³� MON pp;_��y�(�:�L� ^�pϒ~"��qa\EF��ŭ���CL_L�P'�J�İEYLO�GGIN�pu��F���$LANGUAGE �F�abyD <�qL�G�qr�y�a ����xu �e�����P���'0������;��cMCH ;���
��(UTg1:\���� �� �������!�3�E�\�i�{��(���lL�N_DISP �sP�ئ�����OCl4b�RDz�S�A@��OGBOOK tM�d��>A���k�X�܏����������<O�Y���	>F	�Q������N`���O�_BUFF 1-u�me2kE� j�FB�iG�� G>P}t�� ����///C/���~DCS w<�{�=���G���/�/�/�/Z$I�O 1x�{ ğ3D��?*?<?N? b?r?�?�?�?�?�?�? �?OO&O:OJO\OnO@�O�O�O�O�O�%E�PTM�dh�#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogopyo�o-��BSEV������FTYP��_�o�m��RS�h���|��FL 2y=����/��������(TP�����b'�NGN�AM�6%.�V$UP�S��GIh������f�_LOADPR�OG %��%	�T_ARCWEL������MAXUALRM'��A5�̀l�'_PRh��� E�	ˀC��zM����x���,�P 2{�W ت	�aڀ	�|�f4��~��� �������(Ο���3� �(�i�T���x���ï ���ү�� �A�,� e�P�����~������ ƿؿ��=�(�a�s� VϗςϻϞϰ����� � �9�K�.�o�Zߓ� v߈��ߴ������#� �G�2�k�N�`��� ����������
�C� &�8�y�d���������������ćDBG?DEF |$�:!�"�$6 _LDXD�ISAQ�#��#ME�MO_APK�E {?$�
 H �������"ˀISC 1}
$�%��oy�M�����QE_MSTR ~�m~%SCD 1���T/�x/c/�/�/ �/�/�/�/�/??>? )?b?M?r?�?�?�?�? �?�?O�?(OO%O^O IO�OmO�O�O�O�O�O  _�O$__H_3_l_W_ �_{_�_�_�_�_�_o �_2ooBohoSo�owo �o�o�o�o�o�o�o. R=va��� ������<�'��`��MJPTCF/G 1�+]�%������MIR 1e�%Ԁp�@T��q���T�< G ?��%�� t�7�q��i����� ��������1�C�֟ ��j�L�V�x���P��� ��ί��0�T�E � q����8��������� 򿐿���� �B�p� R��ϵ���Z�|���п ����6���>�l�R�d� �߈ߖ����ߌߞ��� 2���@�z�`��� ���������+�=��� �����X�b�t����� ��������*��o �6������� ��
@nP ���Xz��� �4/�,/j/P/b/�/h�/���K������  �/��LTA�RM_�"�̅�� �"����6?>4��METPU  T�����%��NDSP_ADCOLX5�� c>CMNTy? �l5MST ���-�?���!�?�4l5P�OSCF�7�>PgRPM�?�9STw0�1���4܁<#�
gA[�gEwO�GcO�O �O�O�O�O�O_�O_ G_)_;_}___q_�_�_�_�_�Ql1SING_CHK  |?�$MODAQ3����#5veE{�~&bDEV 	���	MC:WlHS�IZEX0�-�#eT�ASK %��%�$1234567�89 �o�e!gTRuI����� l̅%&�O2}��F�cYP�a��9d"c�EM_INF 1��7;a`)�AT&FV0E0�X�})�qE0V�1&A3&B1&�D2&S0&C1�S0=�})ATZ�#�
�H'�O��qCw��A���b�ˏ���� �&��� ����3���ۏȟڟ ������"�4��X�� ���A�S�e�֯៛� �C�0����f�!��� q�����s�俗����� ͯ>��bϙ�sϘ�K� ��w��������ɿۿ L����#ϔߦ�Y��� ��ߩ߳�$���H�/� l�~�1ߢ�U�g�yߋ� ��� �2�i�V�	�z��5����������.ON�ITOR�0G ?�kk   	EOXEC1�22345�`U789 ���(�4� @�L�X�d�Pp�|�2�2�U2�2�2�2�U2�2�2�2��3�3�3(#aR�_GRP_SV �1��{ (�Q��4���Ҿ��~?܉E?��\���+��Ʈa_Ds�n�IO/N_DB-`�1m�1_  �� �Fh�"$ �++��0LFh��N �82)Fi-ud1}e�/�/��/1PL_NAM�E !�e� ��!Defaul�t Person�ality (from FD)b"�P0RR2� 1��L68L@P<�!?`
 d�2-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO@_OqO�O�O�Of#2)? �O�O�O__,_>_P_b_t_f"<�O�_�_�_ �_�_�_
oo.o@oRo�dotl�" �_�n
�o�of$P�o�o  $6HZl~�� ������o�o2� D�V�h�z������� ԏ���
��.�@�� !�v���������П� ����*�<�N�`�r�Ą���e����ïխf"d������� �(�6����� �m���8j���V� ���� ��Ŀֿ�����:Ϸ��]�m�f"��	`ি�ϲ��σ�:��oAb)�����c'? A�  /�	2�3��)X ����E ���X, @D��  t�?�z�n�?xf |�f!AI�tռj��;�	l��	� � � �h�Y �!0���� �� x � � ���ҷK_K �}K7X�K���J��?J�+Ƀ�%��ԯC��@�6@�
��\��(E@�S�����.��=�N��������T;�f�a������$��*  ´�  �1�>��B���z�w����<� 
��� ��!/���1��yD�  ��  �  �
`�#H �l����-�	'� � ���I� �  ��0�&�:�È~��È=�����0�@����%�f���f�(�2�+�a!v  '�Y���@!�p@����@��@��@��C���C� �� C���C��C��f ��A��������9"T�Bb $/��Lf!Dz��o�� ~���������A� �кD�  �X ,f �?�ff0G�*/</� }�q/ă+1�8~`�/�*>�#��$��(�(~`�%P�(������>�$����W�<�	<�S�;�9<���<#*o<c��M,@�K;�|��f��",�?f7ff? ?&�0T��@�.�2�J<?N\��55	��1 ��(�|��?z��?j7�� [/0OOTO?OxOcO�O��O�O�O�O�O{h�5F���O2_�OV_�?w_ �9I_�_E_�_�_�_�_ oooLo7opo[o�o o�o�oU�o�o��m_ 3�_Z�o~���FO*��& Q/�wl�� q
�m.��+�d�V�B��Aa0��5uCP��L�č?��`��#��Y�/Ӄ�6�B]�D��C!C3� z����������@I�l�����A��A��P�A �R?�1�>�-8������ÍO\����Q�߸�#�
؞����AиRA����C;���Q�섟"\)C�0���qBo�
=��Q�����8�Hp��G�� H�0�H���E1� C��&�Hy��I���H��%F��� E,�s�]�i��EI��@H����H��E# D�7�د� կ���2��V�A�z� e�w�����Կ����� ��@�R�=�v�aϚ� �Ͼϩ��������� <�'�`�K߄�oߨߺ� ���������&��J� 5�G��k������ �����"��F�1�j� U���y����������� ��0T?x� u�������P�(�3�(��	4���<��̷�t�Ӂ3�� ���ʭx��Ӂ� &n��
/4�f4y��$-$)d/R/�/v/�/��,ՅPD2P�.�a �o?Z?=?(?a?L<?g?n?�?�?�?�?�??  �����?�? +OOOO:OsO?�o�O�O�O�L7�O�O_�O0 _F_4_JQ�L_^_��_�_�_�_�_�Z  92jOo  B��}�J��Cq���Ӏ@�� RoӀMqko}o�o^o�oҌo�o�o/TAӄ�TӀӀ��aӀ؎
  I������� �)�;�M�_�q�����sq ���1���"�$MSKCF�MAP  $%?� �Vsq�oq莼�ONREL7  �%Ӂ�P���EXCFENBb�
у���FNy��'��JOGOVLKIM�d��d��WKEY�q�z�_PAN��������RUNa���SFSPDTY� '�����SIGN��TO1MOTc�����_CE_GRP [1�$%Ӄ\dO h�\O�����T��ɯ�� ���#�گG���<� }�4�����j�׿���� �Ŀ1��*�g�ϋ� �τ���x����������f��QZ_EDI�T�͇��TCOM_CFG 1�ɍ�~vv߈ߚ�
V�_/ARC_"��%P��T_MN_MOD�E��0�UAP�_CPL��4�NO�CHECK ?ɋ �%�3� E�W�i�{������ ��������/�A���NO_WAIT_�L�K�6�NT^��ɋu|��_ERR�@�2�ɉ�Q�  ��������4�F��MO����|�t5�!�������"�B�o�-B�^����e�<���?�l�Knp����PAR�AM��ɋ��/�2t8�_^ �=�P345678901x��s� ���//�9/K/'+t7�}/�,"�/~��ODRDSP����0�OFFSET�_CARA���&DsIS�/�#S_A���ARK�L�OPE?N_FILE0h����Lִ�OPTIO�N_IO����m0M_PRG %Ɋ�%$*�?�>I3WO�50�F�0� �5���2��0@9�'A	 ���C쯆�#�� RG_DSBL  Ʌ��v|rO�!RIE�NTTO��!C�mpҁ,a� UT__SIM_Du7Ђ���� V� LCT ���H��4���I�%<y��A_PEX��?nTRAT�� d0��T� UP ��N�pK��i_{_Xr�fS`�gq�2m�}]��$�2?��L6�8L@P�C
 d�/�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J\��2�_���� ���
��.��{ X�j�|�������ď֏ �������H�X��PX�~��"Pk����� ̟ޟ���&�8�J� \�n������������� ����"�4�F�X�j� |�������Ŀֿ��� ɯۯ0�B�T�f�xϊ� �Ϯ�����������`,�>���E�}���SI�߿ޤ��� ��b�bݢ/3��W�
�@L�v�l�~��� ������J�Q�'�)L�	``�Z�l�~���:�o�A������|��KA�  ����T�POOP1��[�v��T�H��E=D�X, @D��  2��,?��D4429�h;��	l�	@�� � �h�_`� ��� � x � �� ��JH��H2�-HL���H�lH�WG���=�3Ho�X�JC��@p�@�ז@�P1��j�0@�S �>PP%ICUB��<��K��@���a�y�  ��  �  +� #�0�*&��H/�	'� �� f"I� ��  ����=���͊/�+�@��/� �>A�/M+>B����N�@4?  �'x0L4�0C�@C��� CC�C��Y?k?D�  ��A�!���������B�@�1�����!
ENz�-O�QO<O�aO�O^/p(�1�E�Sȇ �<��1�P.  ? �?�ff��O�O�O 7�/_A[sAq8�W_eZ>�'� �FjJ(��UP �X�I����#�T[���<�	<�S�;�9<���<#*o<�1�5�\@�	k:���#�R��?ff�f?� ?&D`�@��.Vb�J<?N\�be:��2?aK jI:�o8�o(g~_ �o�o�o6!ZE ~�{����� ��o�o�o�h���� w�����ԏ��я
��� .��R�=�v�a�?�� o�e+��O����<�0N�`�r�Z���@_��l� /�ȯ+��ׯ�"����A`>��?��C�s�
�П��?�ء����̿n	[�/X���B��D90CC�ޚ���x����^�@I�*�����A��A���PA �R?�1>�-�������ÍO\����Q�����#�
������AиR�A���C;����Q�B��0\�)C0����qBo
=��Q�������Hp���G� H��0�H��E1� C���Hy���I��H���%F�� E,��1߯i�EI���@H���H���E# D� ���ߨߓ��߷����� ���8�#�5�n�Y�� }������������ 4��X�C�|�g����� ����������	B -fxc���� ���>)b M�q����� /�(//L/7/p/[/ m/�/�/�/�/�/�/? �/6?H?3?l?W?�?{?��?�?�?�?�?O��(Ζ�3�([��T��<BE�5�̷�2ODOX�3���^OpO~B��ʭ�O�OX�� �&n�O�O4�f4yϱ�M�I"__�F_4_j_X\��PbP�^�����_O�_�_�_o
l?%o,oeoPo�uo�o�o  ���ʞo�o�o�o�o1@�_��dR�v|7�����������
��R�@�v�d���Ψ�  2(я  QBG�;�G�C/�D�X�@K��"�4�F�X�j�{���������ɟP۟���X���X��X���X���
 �W�i�{����� ��ïկ�����/��A���1� ���K1���"�$PAR�AM_MENU �?�E��  MN�UTOOLNUM�[1]݆��F�~�����AWE�PCR��.$INCH_RATE���SHELL_C�FG.$JOB_�BAS߰ W�VWPR.$CENTER_RI�������AZIMUT�H OPTB�����ELEVATI_ON TC�����DW�TYPE �SN�ARCLI�NK_AT �ST�ATUSǳ]�__�VALU߱̰L�EP��.$WP_ �����U�̢ϴ����� �����7�2�D�V���z�SSREL_IOD  �E�Q����USE_PROG %��%{��ߏ�CCRT�ԶQ�����_HOST !F��!��5���T�P��Q��*�S����_TIMEOU��  z�GDE�BUG�Љ���GI�NP_FLMSK̶���TR����PG�d�  ����$�C�H����Q��� z�tߪ��������� (:c^p�� ����� ; 6HZ�~��� ���// /2/[/���WORD ?	���
 	RS��CPNn�BgMAIW��#SU&��#TEt�CSTsYL COL0e�W(�/W�TRACE�CTL 1��E��� �P |��6DT Q��E�D0!0D � ��S��Q�Q6�[<��Qy01�q?�?�?�? Q5�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c�u��������� Ϗ����)�;�M�0_�q�S36LEW���v5��3  �6?_UP �<;b�s����� ���&�0�M$a��R�\0�R�  ��)_�DEFSPD ��2��  ��z�INؐTRL' ���a�8!�h��PE_CONFI:ܐ�7���M!]b,LIDٓ����	ĨGRP 1��9 lM!A>ff��\��
=D�  D_Z� D
�@�
�M d!�?�O�������H�"�$�i�G ´����m�B�� ̱�������̿��&�B34�$��]�o�Y� <<j ��tϭ�pϪ������ �ό��O��_߅�p�"�z�ӳ�M 
���� �������5� �Y�D� }�h��������������*�)<�
V�7.10beta�1�� A�k=�\�B
��(�Y��?&ffp�>.�{X�
������X�B!념�A{�33A�&�(�h� @-�����������pM"��3EWM$�ғ�KNOW_M�  0��ȤSVw �:�%��������IM"G��M��=�(�	������.�* �����M#�)�Y�@)���M %X .ѐȡMR�=��$����f/x+��S�T�1 1�<9^ 4�()�o��/ �/�/
?�/?!?S?E? W?�?{?�?�?�?�?O �?�?>OO/OtOSOeO�wO�'2�,��/���#<�O�O� 3�O�O�O�O�'4_-_?_Q_��'5n_�_�_�_�'6 �_�_�_�_�'7o&o8oJo�'8goyo�o�on�'MAD�� ȕ��EOVLD  ����P}�$PAR?NUM  �+?�Q�#SCHy �ȕ
�wlq�y��uU�PDl=u���E_CMP_u����_��'ݥ%�ER_CHK3�ۣ �G�0��B�RSA �ȡ_M�Op����_���E__RES_G� ���
��p�"��F�9�j� ]�o�����ğ���۟@����o��@��� 1��PN�m�r��mP ��������P̯�� �`�*�/��f`J� i�n�惹`������悏V 1���ށ��@]s8��THR_INRA �q]م�d�MASS)� �Z=�MN(�[�MO�N_QUEUE C������!ބN*�Un�NkƔȫ��END��Ώ��EX1E�����pBE����>��OPTIO��׋���PROGRAM7 %��%�������TASK_I�t �OCFG ᯎπ�ߵ�DAT�Ax����G2 �$�6�H�Z�l��� ����������� ��2���INFOx�혝���������� ������	-?Q cu������h�N�Z��� �l���pK_����ٴz�5G��2�D� X,		x��=����@	���$� �����0_EDIT ��������WE�RFL��Ó#RG�ADJ ��A	Л@R$?�]%0�5&���?���'�?���A<��z�%�o�/)(/s#�2�'"	H��l��!?8��Aٴ�t$26�*A0/C2 **:@L2�??Q3m=���2F�5��+1�9��/ �?y=�=�?�?�?�? �?KO�?O5O+O=O�O aOsO�O�O�O#_�O�O ___�_9_K_y_o_ �_�_�_�_�_�_�_go o#oQoGoYo�o}o�o �o�o�o?�o�o) 1�Ug���� ����	���-�?� m�c�u����ُϏ �[���E�;�M�ǟ q���������3�ݟ� ��%���I�[���� �����ǯ������	�ߖ�𰄿����39 ߿53��ϧ�0�B�o'PREF �*�00
5%IOR�ITY:���9!MPDSP8�'*z���UT��34&ODU[CT���E�v�&OG_TG$ ������TOENT� 1�� (!AF_INE���Y�J�!tcp|dߌ�!ud{�~��!icm�߬�.��XYx#���1)� Y1�*�0��S�6�B�� f������������!�3��W�>�{���*��x#�)P�/������Y7/c<��4�4��(�.A�",  �u�(}� ��+%�^Ŀf�x��,9!PORT_N�UM��0��9!_CARTRE�P% �aSKST�A�� 4LGS6V�����#0�Unothin�g����L�]T?EMP �����T��_a_seiban�,/�</ b/M/�/q/�/�/�/�/ �/�/�/(??L?7?p? [?�??�?�?�?�?�? O�?6O!OZOEOWO�O {O�O�O�O�O�O�O_ 2__V_A_z_e_�_�_��_�_�_�_�_o�VOERSI����M`� disab�led'oSAVE� ���	26�70H782J�o�o!$�o�o���oC 	x��V��.�eKt���J�Ac|�o���mb_�W 1����`*��p�!�4�F��W�UR?GE_ENBЪ�l(���WFr�DO�Ƅ�+�WRГ���W�RUP_DELA�Y �,��R_?HOT %{����#���R_NORMAL����W�&�SEMI6�\���U�_QSKIP���#�xo��	o��(� ��Y�G�}�����g� ů��կ�����C� 1�g�y���Q������� ���	�Ͽ-��=�c� uχ�Mϫϙ������� ���)��M�_�q����$RBTIF���0RCVTMOU�E����DC�R�Ǿ� ����6uC^�)C7��@����@�n�6����띶��^���R�����-���j����H�3�<�	<�S�;�9<���<#*o<��M�Q 7���y��������/��A�S�e�w������R�DIO_TYPE�  ����EFPOS1 1�ui� xA
-���G 2k�o�*�N� ���1�Ug N���n� �/�/Q/�u// �/4/�/�/j/|/�/? ?;?�/_?�/�??�? �?T?�?x?O�?%O7O��?�?OOjO�O��O_S2 1�ԋ�ZO�O_�O6_�O��3 1��O�O�O,_�_��_�_L_S4 1� c_u_�_�_?o*oco�_S5 1��_
oo�Vo�o�o�ovoS6 1͍o�o�o�oiT|�S7 1�"�4F���"��S8 1Ϸ����~���5�SMAS/K 1���  �� �ՇXNO���)�x=�����MOTE���=�Z�_CFG ��a���)���PL_RANG]��ߛ�OWER �%��ΐ��SM_DRYPRG %%��%^��ԕTART� �ƞ�UME_PRO���p�=��_EXEC_EN�B  ���GS�PDI������Ѣ�T3DB����RMϯ���IA_OPTIO�N������U�MTE_݀T��_���*�fz��9���C�ˀ�����������OBOT_ISOKLC"�����ֵNAME %��_���OB_OR�D_NUM ?�Ƙ��H7�82  ˄h�@�h�$�hʬ�h�>�P?C_TIME�םٽx��S232z�1�����LTE�ACH PENDcAN��v�A�~��]�H@Maint�enance C�ons˂��ˆ"��DDNo Use~�E��i�{ߍߟ�8�ߵ���NPO#����A�!���CH_�LL��U���	�3���!UD1:�Y� �R܀VAIL�I����U�SRW  %������R_INTVAL����������V_DATA_GRP 2�%���X�D��P��W���{� f�%������������� ��$&8n\ ������� �4"XF|j� ������// B/0/R/x/f/�/�/�/ �/�/�/�/�/?>?,? b?P?�?t?�?�?�?�? �?O�?(OOLO:O\O ^OpO�O�O�O�O�O�O�_ _"_H_6_l_U���$SAF_DO_PULS��V���X���Q�PCAN������SC���(�����ˀq�����x�C�C��˂  p�o0oBoTofoxoo��o�o�o�o�o�o������be�!r �d�t:ql�(s�� @��fx��~Ny�� D�t�_ @�T�������T D�� *�S�e�w��������� я�����+�=�O��a�s�����`u2���ǟі��C�^��;�o2����p����
�t���Di���aC��  � ���Cђa x��Qa�s��������� ͯ߯���'�9�K� ]�o���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ�����������1�2��aZ�l� ~ߐߢߴ�������9� u�(�:�L�^�p��@�������2�0� D��N�	��-�?�Q� c�u������������� ��);M_q ������� %7I[m� ����D��/!/ 3/E/W/i/{/�/�/
� �/�/�/�/??/?A? S?������r�?�?�? �?�?�?�?O#O5OGO YOgIzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_�oo*o<oNo`o5�� ��9�ko�o�o�o�o�o &8J\n� ����pj�o�\�2���S�����	12345�678+�h!B�!ܺ�4���`��|�������ď ֏������o5�G� Y�k�}�������şן �����1�C�U�f� $���������ѯ��� ��+�=�O�a�s��� ����h�z�߿��� '�9�K�]�oρϓϥ� ���������Ͼ�#�5� G�Y�k�}ߏߡ߳��� ��������1�C�U� �y���������� ��	��-�?�Q�c�u� ������j������� );M_q�� �������% 7I[m��� ����/!/3/E/ W/{/�/�/�/�/�/ �/�/??/?A?S?e? w?�?�?�?�sm��?��?q/OO*OF��Cz  Bpqj �  ��h2�b�m�} ph
�G_�  	��r2�?`�O�O�O�Ook>�_D	lo�<��OB_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o'_�o�o�o�o (:L^p��� ���� ��$�>I�SB�1�AiB<S���$SCR_GR�P 1��8�� � � }�SA dE�	 ����������1B����SG��ۏɏ�:Mi�s@��D^@D/^�E��� \AR�C Mate 1�00iD/145�0ҁAM�ҁ�MD45 678�SC
12345��9��ӅE����KyBד_��SF�߃�@ S��Ó��Ӂ�	yJ�6�H�Z�l�~�SD���H������ ���Əǯ���Ά�oSAگC�֯g�N���v�B�M@Ʋ���ɴr��A^@ؿ  @S@�𵬁@��� ?PŬ�HM@)�ۺ��F@ F�`S� [�~��jϣώϳ��� ������!ߤ�� �L�07�I�[�m�B�{�� �߬�����	����?� *�c�N��r��_�� )������dG�@���0�SB�@P7H��_�!�@�p�M@�������߃�?���SDA�������$�� QƒSA 3E��!ht�U (� ������� �$SF_�E�L_DEFAUL�T  ����S@@HO�TSTRL#^�E�MIPOWERFL  BEX?�oWFDOM ��RVENT 1������w L�!DUM_EI�P.���j!AF_INEL/SDO!FT�@./rd/!���/ �S/��/!RPC_M'AIN�/�(��/�/N�#VIS�/�)��/�H?!TP;0PU�??�d7?�?!
P�MON_PROX	Y�?�e�?�?[2�?��f�?,O!RD�M_SRV-O�gOxO!R���O�YhgO�O!
� M�?��i�O_!RL�SYNC_��8|�O\_!ROS��\�4K_�_!
C}E]0MTCOM�_��k�_�_!	�RC'ONS�_�l�_@o�!�RWASRCdGO�m/o�o!�R'USB�o�n{o�o w/�o;C�o�o%J�n5�Y�:RV�ICE_KL ?�%� (%S?VCPRG1���"�u2�
��p3-�2�"�p4U�Z��p5}���"�p6�����p7͏ҏ��p����9�"� �t�OJ��q�r��q� ���qG��qo���q ����q��:��q�b� �q����q7����`� گ�������*�� ؟R�� �z��(��� �P�ʿ�x����� ��ȯB�D����r �p��p����<����� ���	�B�-�f�Qߊ� �߇��߫�������� ,��>�b�M��q�� ����������(�� L�7�p�[�������� ��������6!Z lW�{�������2V�z_�DEV ���MC:��T4���pGRP �2�����pbx� 	� 
 ,�^����/� &///\/C/�/g/�/ �/�/�/�/�/?�/4? ?X?j?��?E?�?�? �?�?�?OOOBO)O fOMO_O�O�O�O�O�O �O�O_q?_P__t_ [_�_�_�_�_�_�_o �_(ooLo^oEo�oio �o�o�o�o3_ �o 6ZAS�w� ������2�D� +�h�O������oy� ���ߏ��@�R�9� v�]�������П���� ۟�*��N���C��� ;�����̯ޯů�� &�8��\�C�����y� ����ڿ��ӿ�g�4� F�-�j�Qώ�uχ��� ���������B�)� f�x�_ߜ߃�����)� �߭��,��P�7�t� ��m��������� ��(��L�^�E����� w���o����� �� 6ZlS�w� �����D.��d Ԗ�	2{�f�����O%���/����� 4!�4%D/R'</r/`/ �/�/�/�)/�/0)�/ ??>?,?N?P?b?�? �/�?�/�?�?�?OO :O(OJO�?�?�O�?pO �O�O�O�O_ _6_xO ]_�O&_�_"_�_�_�_ �_�_oP_5ot_�_ho Vo�ozo�o�o�o�o(o Lo�o@.dR� v�� �$�� �<�*�`�N������ ��t���p�ޏ��8� &�\�����L����� Ɵȟڟ���4�v�[� ��$���|�����¯į ֯�N�3�r���f�T� ��x��������:�� J��>�,�b�Pφ�t� �����Ϛ�ߖ�� :�(�^�L߂��ϩ��� r����� ����6�$� Z�߁���J����� �������2�t�Y��� "���z����������� :�1��
��R� v����6� *:<N�r� ���/�&// 6/8/J/�/��/�p/ �/�/�/�/"??2?�/ �/?�/X?�?�?�?�? �?�?O`?EO�?OxO 
O�O�O�O�O�O�O8O _\O�OP_>_t_b_�_ �_�_�__�_4_�_(o oLo:opo^o�o�o�_ �oo�o �o$H 6l�o��\~X ��� ��D��k� �4����������� ��^�C����v�d� ������������6�� Z��N�<�r�`����� ����"��2�̯&�� J�8�n�\���ԯ���� ���~���"��F�4� jϬ���пZ��ϲ��� ������B߄�iߨ� 2ߜߊ��߮������� �\�A��
�t�b�� ������"����� ����:�p�^������� ������� "$ 6lZ������� ��� 2h ���X���� 
/�/p�g/�@/ �/�/�/�/�/�/?H/ -?l/�/`?�/p?�?�? �?�?�? ?OD?�?8O &O\OJOlO�O�O�O�? �OO�O_�O4_"_X_ F_h_�_�O�_�O~_�_ �_o�_0ooTo�_{o �oDofo@o�o�o�o �o,noS�o�t ������F+� j�^�L���p����� ��܏��B�̏6�$� Z�H�~�l����
�۟ ������2� �V�D� z�������j�ԯf�� 
���.��R���y��� B�����п������ *�l�Qϐ�τ�rϨ� ���Ϻ����D�)�h� ��\�J߀�nߤߒ��� 
������ߴ�"�X� F�|�j�������� ����
���T�B�x� �����h��������� P��w��@ ������X ~O�(�p�� ���0/T�H/ �X/~/l/�/�/�// �/,/�/ ??D?2?T? z?h?�?�/�??�?�? �?O
O@O.OPOvO�? �O�?fO�O�O�O�O_ _<_~Oc_u_,_N_(_ �_�_�_�_�_oV_;o z_ono\o~o�o�o�o �o�o.oRo�oF4 jXz|��� *���B�0�f�T� v���Ï������ ��>�,�b�����ȏ R���N�̟����� :�|�a���*������� ��ȯ�ܯ�T�9�x� �l�Z���~�����Ŀ �,��P�ڿD�2�h� Vό�zϰ�����Ϡ� �Ϝ�
�@�.�d�R߈� �ϯ���x��������� �<�*�`�߇���P� ������������8� z�_���(��������� ������@�f�7v� jX�|��� �<�0�@fT �x����/ �,//</b/P/�/� �/�v/�/�/?�/(? ?8?^?�/�?�/N?�? �?�?�? O�?$Of?KO ]OO6OO~O�O�O�O �O�O>O#_bO�OV_D_ f_h_z_�_�_�__�_ :_�_.ooRo@obodo vo�o�_�oo�o�o *N<^�o�o� �o�����&�� J��q��:���6��� ڏȏ���"�d�I��� �|�j�������֟ğ ��<�!�`��T�B�x� f�������ү���8� ¯,��P�>�t�b��� گ��ѿ�������(� �L�:�pϲ���ֿ`� �ϸ�������$��H� ��o߮�8ߢߐ��ߴ� ������ �b�G��� z�h��������(� N��^���R�@�v�d� ������ ���$��� ��(N<r`��� ������$ J8n���^� ���/� /F/� m/�6/�/�/�/�/�/ �/?N/3?E?�/?�/ f?�?�?�?�?�?&?O�J?L1�$SERV�_MAIL  �T5J@�0HOUT�PUT?H}0HRV 2��6;  M@ (�1O��O4DTOP10 �2�I d  P?�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o��������5�EYP�E`LNEFZN_C�FG ��5�MCL4oB�GRP� 2�%�� ,�B   Ae�L1D�;� Bf�� � B4L3RB{21�FHELL�C��5��@�O<�|ΏK%RSRݏ ޏ��)��M�8�q�\� ������˟���ڟ����7�I�[��  �+�[�����i��� L0��ŢơL8
q�2L0d��������HK 1瞋 ˯@�J�D�n����� ����߿ڿ���'�"π4�F�o�j�|ώϊ�OMM 螏�Ϗ��FTOV_ENB�?D�A��OW_R�EG_UI��2BIMIOFWDL������h�3�WAIT�����oE^�Z@�܇DX�TIM������VA>@i�3�_�UNIT�����L]C�TRY���4@MON_AL�IAS ?e���@heOM�_�q�� J;����������  �2�D�V��z����� ����m�����
. ��Rdv�3�� ����*<N `�����w �//&/8/�\/n/ �/�/=/�/�/�/�/�/ �/"?4?F?X?j??�? �?�?�?�?�?�?OO 0O�?AOfOxO�O�OGO �O�O�O�O_�O,_>_ P_b_t__�_�_�_�_ �_�_oo(o:o�_^o po�o�o�oQo�o�o�o  �o6HZl~ )�������  �2�D��h�z����� ��[�ԏ���
��Ǐ @�R�d�v���3����� П⟍���*�<�N� ��r���������e�ޯ ���&�ѯJ�\�n� ��+�����ȿڿ쿗� �"�4�F�X��|ώ� �ϲ���o������� 0���T�f�xߊ�5߮� �������ߡ��,�>��P�b���$SMO�N_DEFPRO�G &������ &�*SYSTEM*�i����<�{�RECALL �?}�� ( ��}3xcopy �fr:\*.* �virt:\tm�pback��=>�192.168.�56.1:13648 � �2�D��}4��a������������ }8��s�:orderfil.datv������/AS}/��mdb:s���� �`���z���.@ Re������� ����~�*/</N/a s/��/�/�/�r �&?8?J?]o ? ��?�?�?��v// "O4OFOY/k/O�/�O �O�O�/�/|??�O0_ B_�Og?�O
__�_�_ �_�?�?�O�O,o>oPo cO�_�Oo�o�o�o�O t_�__(:L__�o �_����_�_xo o$�6�H�[omo��o ����Ə�o�o~ � 2�D�Wi������ U�������.�@� R�e� ��������Я �v����*�<�N�a� ��������̿ߟ� z��&�8�J�]�o�
� ���϶���ۯ��� "�4�F�Y�k��Ϗ��� ����׿����ߟ�0� B���g������� ����x߅��,�>�P� c�����ߪ������� ��|��(:L_�s� ��������� �$6H[�m���� �������t� / 2/D/Wi/�/�/��/U.�$SNPX�_ASG 2������!��  0�%���/?  ?��&PARAM ��%{�! �		;�P���o4��� OFT_KB_CFG  ���%�#OPIN_S_IM  �+j2��?�?�?�3� RV�NORDY_DO�  t5�5BQSTP_DSB�>�j2HO�+SR }��) � &n:�O��&TOP_?ON_ERRO�F�PTN �%��@�C�BRI?NG_PRM�O#B�VCNT_GP �2��%l1 0x 	DO?_�-_f_Q_�_��'VDPRP 1	�C9m0{Q�1m_�_ �_�_�_o4o1oCoUo goyo�o�o�o�o�o�o �o	-?Qcu �������� �)�;�M�_������� ����ˏݏ���%� L�I�[�m�������� ǟٟ���!�3�E� W�i�{�������دկ �����/�A�S�e� w���������ѿ��� ��+�=�d�a�sυ� �ϩϻ��������*� '�9�K�]�o߁ߓߥ� �����������#�5� G�Y�k�}������ ��������1�C�U� |�y������������� ��	B?Qcu����RPRG_CoOUNT�6��BN�	ENB�O�M���4�_UPD 1}�nKT  
� �ASe���� ����//+/=/ f/a/s/�/�/�/�/�/ �/�/??>?9?K?]? �?�?�?�?�?�?�?�? OO#O5O^OYOkO}O �O�O�O�O�O�O�O_ 6_1_C_U_~_y_�_�_ �_�_�_�_o	oo-o VoQocouo�o�o�o�o �o�o�o.);M vq������ ���%�N�I�[�m� ��������ޏُ돷�_INFO 1�,/ �� �R��=�v�a������!�������"��B�o-B�^������YS�DEBUG� 0����d��SP_PwASS�B?�LOG �/]9  ������  ���UD1:\���_MPC$�/�����/[�Я /��SAV �'�����G�_���f�SV�ԛTEM_TIM�E 1�'�:k 0� ����ү�r�4�SKMEM � /�G� � ��%s���Ͽ��� @����������M"��P׿A��A�;��D�V���n�������Ϧϸ���r^��E�� W�������+�=�O�a�s� �ߗߩ߻����������{�9�K�]�o�� ������������� #�5�G�Y�k�}����T1SVGUNS�*�'���A�SK_OPTIO�N� /���_�DI����BC2_GRP 2�/��Q�%��@5�C��:��BCCFG 3�� ����`������ ��!E0iT �x�����/ �///?/e/P/�/t/ �/�/�/�/�/?��, !?�/T?f?�/C?�?�? �?�?�?׮O���0O 2O OVODOzOhO�O�O �O�O�O�O�O_
_@_ ._d_R_t_�_�_�_�_ �_�_o�_oo*o`o Fh10to�o�o�o�oFo �o�o�o"FXj 8�|����� ��0��T�B�x�f� ������ҏ������ �>�,�N�P�b����� ��roԟ���(��� L�:�\���p�����ʯ ���ܯ� �6�$�F� H�Z���~�����ؿƿ ����2� �V�D�z� hϞόϮϰ������� �ҟ4�F�d�v߈�� �ߚ߼�������*� ��N�<�r�`���� ���������8�&� \�J�l����������� ������"XF |2ߔ����f �B0fx� X������/ //P/>/t/b/�/�/ �/�/�/�/�/??:? (?^?L?n?p?�?�?�? �?��?O$O6OHO�? lOZO|O�O�O�O�O�O �O_�O2_ _V_D_f_ h_z_�_�_�_�_�_�_ o
o,oRo@ovodo�o �o�o�o�o�o�o <�?Tf���& �����&�8�J� �n�\���������Ə ȏڏ���4�"�X�F� |�j�������֟ğ�� ���.�0�B�x�f� ��R��Ư������ ,��<�b�P���p����A��*SYST�EM*��V9.0�055 ��1/3�1/2017 �A v  ��K��TBCSG_G�RP_T   �\ $ENAB�LE�$APP�RC_SCL �  
$OPE}N�CLOSE�S_MINF2'��ACC��PAR�AM� ���M�C_MAX_TR�Q�$d�_MG�Nk�C�AVw�SwTALw�BRKw��NOLDw�SHO�RTMO_LIMȺʧ�h�J����PLQ1��6���3��4��U5��6��7��8k������� )$D�E�E��T��b�PATH^�w�m�~w�_RATIOk��s�T� 2 	/$CNT�A������m�INX�_UC�A���CAT_�UM��YC_ID� 	����_E�����6������PA�YLOA��J2L�_UPR_ANG6�LWA�?�3�O�x��R_F2LSHRTv�LOD���}��������ACRL_S��ؽ���+�k�HVA��$Hx���FLkEX�B�J2�w P�B_F��{$��_FTM���&��$RES�ERV�>�;������� :$��LEN.�z�;�DE|���;�Yғؔ����SLOW_AX�I��$F1��I���2��1������MOVE_TIM��_INERTI���
�	$DTOR�QUEX�3��#I>��ACEMN��%(E�%Ep	V��d�pA�R�TCV���Rt����
��T"@�RJ���	�M��,��J�_MOD�����S dRy�2��	PpE���\��X��AW�gQJ�K@��K��VKv�VK�JJ0����JJ�JJ�AmA��AA�AA%f�AA �t�N1��N �d�#��E_N�U��A�JCFG�� � $GoROUPc�SK��_B_CON�C���B_REQUIR�E���BU��UP�DATT�E�L}  �%� �$TJ��� JEΤ�CTR��
TN� F�&�'HAND�_VB��OPn� $oF2x��3�m�COMP_S�W�#B�R�� '$$Ma�e�R�Î8����<� �5�¼6A_�.�h�D�<q�A��A���A��A���0��D���D��D��P��GR�ǂAST�ǂA���AN��DY���x� �4�5A���s��s��2�B��R����P ����� �)�2�;�s�h�� �0i�\� 7�U6��QOASYM��
�T�¡��мݎ���_SH�"�������TU8����%�7�J>���P�ppcfio�_VI83��h6þ`V_UN!I���d�{�JU�b U�b���d���d v����������su�|�� ����T�oHR_T��	N2��q���DI����Op�t@Ңp�#
  
�2I�QAz����q ��S�s � B� �p � � f1M�Ee���pr�QT�pPT&`r a�>����~$�5`C�^�R�T�4`! $DU�MMY1�$P�S_ RF��u$����FLA� �YP_��F�$GLB_T�0�u΅>����1�:1�q �X��'�STf�� SBRv�M21�_VT$SV_�ERa�O(`�,�C)L��Ap O�r�p�GL�`EW� �4 $H�$Y
�2Z�2Ww��x�b3�A���@�Y�U]�� oN��)`$�GI0}$]� �d�W���� L�h���'b}$F'bE^��NEAR_ N��yF�\ TANC���@�JOG���� �e�$JOIN�T�& ��MSET.�  ��E��� S��@̔� ���  Ue?��� LOCK_F�O��m1�pBGLV�3GL��TEST�_XM�j�EMP�=�Ϣ悖�$1UC�\���2� ��B����i0������CE| Ó� $K�AR�M�sTPD�RA`�3�*�VEC�~�D�.�IU���!C{HE��TOOL���i�V��REK�IS�3;���6���AC)HP���v�O��F����29���I�� � @$RAIL__BOXE�� oROBOƤ?��?HOWWAR���<����ROLM��ŀq!��¡!Ӱ��J�O{_F� ! =1�Y���K�6� �R
N�Oo�W���?�C�Y�sZ�OUR������Q�"�!��$PIPǦN]�Ӳࣱ ��V�@�CORGDED����u��p�� O�p  D ̀OBA�#��������̀��'`�!S;YS��ADR�!�p�>�TCH�0 � ,oEN�r#�A���_��d�z!�%P�VWVA� Ǥ 9�]��uPR�EV_RTA$�EDIT��VSHWR�!�&��]q�%�`D(�.Q��6Q?$HEAD8amp4��Ha��KEq�|��CPSPD�JM%P�L�u�Ra �t����\�IРS�"C20NEr��!�'OTICK���QM�Q�f�:�HN��� @�W�~%�_GqP��ʶ$�STY^���LO�5�8���_ t 
��Gj�S%$�Ѳ�=��S�!$�aJp-����pr��P�P��SQU-�x�����aTERCB��"��TS�$ ����']�'-`�b>pOC�6�bPIZ��4������PR�������S��PU�a��_�DO�c�XSN�KN�vAXI��/���UR� p�"찕�"�d]1� _`�4�ET5QP��ЦU��F�W2��A�A�Q��ĳ���!�h�RE4lu��9��:� �6�	�2��7��9� �9�G�G�'F "TIF�R&��4CE o2oDoVd�!�SSCЀ  �h� DS��4���S�P�p"%AT@�2����c⅂ADDR�ESs�B��SHIyF�#�_2CH� ��I�t!�TU��I�1 W�C�USTOV �+TV��I�r UҸ�h6!��P
Ϫ
�s1qV������! \���������,��J�2C�SC��Y�*��2�1�TXSCREE���"�p�TINAO���T4���q66"vP# TI�/���4� .���63��4��RRO�@�3�
��1����UE?�$ �ȍPMѧ�SP�4�RSyM����UNEX_��vA�pS_��+F�S A.IIG�S6C��Bވ4 2#O0UE�rT%�r?�nF��GM�T3pL�a�O�@�6�BBL_��W�o���& ����BO���BLEf"�C밼�"�DRIGH�CB�RDA�\!CKGRo�UTEX$ UQWIDTH�����Ʊ��Jq �UI�>�EY6 ��' d�h��Ѐ���Ӱ��B�ACK�ᡂ�UE��!�FO���WLAB��?(!�I����g$UR��P m^Q�'�H�1 ( 8�wq�_��t"�R(�R�q�����������QO�m!��)��L�PU��@7cR���LUM87cV ERV��U�R_PP�fT*�j CGE�R�a `�)��LP�e_E\���)��g��h!�h���i5*�k6�k7�k8�bZ�@6����4�������SJ�)^QUSR�]�+ <��'�U����#��FO� ��P�RIrm��%q�pTWRIPϱ�PN�p
�t,����p����p/��3 -� -�R\Sp��G  �T/���u!�rOSF��vR 9 �2�so���.f�x� ����h��U�a���/$�6�DC�b���sOSFFŠ��0��L�=O�� 1.9���Z��/9�GU.�P���׃��sQSUB8��H��@SRT��a1���;���OR��N'�RAU� (�T=��Z��VC� Ҕ2G� ɲ��$����y�8񹳬`C��{�D�RIV��@_Vа����Ѐ�D4tMY_UBY3t����� $��19�l0��	����P_S������BM�A$b�DEY_�EX�@�3����_MU.�X�An� @USA8��p[�k0w��xp� �2x�GgPAgCINr�!�RG�� ��������A���SCp�CRE�Rj!o��`�ܽ�S�3 Y�TARGÐP�"��pa�	R�S�4nP0`TQ��	o���REz�SMW��_A��� o���OIq\!An v��EE$pU�෱� \PVa�HK��5����`W�s��0��EA��ɷWOR�Pv��P��MRCV�A6 ���`O��M�PC�#	p����REF�G (����e�s`cM�Xp �^��^�-ˀ�Ƶ��_RCʻ���0S !pf�ϓ��a��D7 ���gPTU0 epԕw�OU�����枃� 2��2� $U00��r�4�5#�^�K SUL6b�5c`CO�0 `6`�]��Ӥ0����@��a��@q��i�L����$���a��@q�|s�?�8| +5#�k� 5#CACH��LOR�&�<�a�A��KQC ��C_LIM-Ig#FRj�Tl�N��$HO�P�*�OCOMM��BO�@���ب �a��VPH��/ ��_����Z�����k���WA{�MP��FAIk�G���;�AD?�p�IMR1E�_���GP@V��� k�ASYNBU=Fk�VRTD����l��&SOLo D_|���WA�P�ETU�O�X�Q����ECCU�VEM٠%�k�VIRC?����|B��_DELA�����p�p�AG��R�c�XYZM@5Cc�W3�qsQ T��P���s��D9�"�QLAS�AP�
�� Gl� :��rX�Sa�7�N�
��VLEXE�;Ȕ3W�ka5!��FL2PIW���FI����F���]�:#
�<_p�
��8t@s\���@ORD|q����##�� =_0Z`T��r�B�OJP6b��VSFE �3> a a0s���c�UR��n�@VSM�u?�rdV�R J� f��"�Ɗ5@�r��qLI�N��@�WN�XSD屎 A��2��K&S]Hd`HOLk�XVR�tB��@T�_OVRk �ZABC�C��"q�-1��Zހ�tD�rD/BGLV��Lϒ�R��P�ZMPCF"�E�0�t2ޑLN~ ��
2d���F Ђ`��ɰ4C�MCM��C��CAgRT_Y1��P_2`? $Jw3q4D��}2�2�7`�5`抲UX|5UXEu��6|�5�4�5�1��1�9�1�6�Z�%gG +�$ �p�AYV D�p Hb�RRM�{q��HETH����PU'�Q�!}P�I � �83�� PEAKf���K_SHI�B��'RV F�G½B� C�@r2g1|�����A�20��I S��DXT/RACE�PVw��B�SPHER'aJ� ,e�THjO|I���$TBCSG� �2 ����Q�����0 
30` �_�_�_�_ �_�_�_�_.ooRodk�wR~S�\d ���a?�Q	 H�CBdo�iC  �B �R�o�h�o�kB���op��o�jdf  AXp?�w {qW�{������@�@0:nT�g� z�E�W���������
���3�	V�3.00�R	mwd45�	*U��M����1�� 8��m���  ��֟,�wQJ2{c�]6�����  �Ue�Q ����E�9şp��p�����	_�ȯ���ׯ� ��4��D�j�U���y� ����ֿ�������0� �T�?�x�cϜχϬ� �Ͻ�������>�P�X�7�j�|�&ߜ��� ������	���-��Q� c�u��B������ �����U%�7��Q�� =�c�Q���u������� ��������)M; q_������ �7%GI[ �������� �//�M/;/]/�/ q/�/�/�/�/�/?? %?�/I?7?m?[?}?�? �?�?�?�?�?�?!OO EO3OiOWOyO�O�O�O �O�O�O_�O__/_ e_S_�_w_�_�_�_�_ �_o�_+ooOo=oso �o//�o�o5/ko�o�o 9'Io]� ��u����� 5�G�Y�k�%���}��� �����׏���1�� U�C�e���y�����ӟ ������	��Q�?� u�c���������ͯ� ���o�oA�S���+� q�������ݿ˿�� %�7�I�[���mϏ� �ϣ����������3� !�W�E�{�iߋߍߟ� ����������A�/� Q�w�e������� �������=�+�a�O� ��s�����e������� ��'K9[]o �������# G5k}��[ �����//C/ 1/g/U/w/y/�/�/�/ �/�/	?�/-??=?c? Q?�?u?�?�?�?�?�? �?�?)OOMO_O��wO �O3OaO�O�O�O�O_ _7_%_G_m__�_O_ �_�_�_�_�_o!o3o Eo�_ioWo�o{o�o�o �o�o�o�o/S Acew���� ����)�O�=�s� a���������ˏ�O 	��-�׏]�K���o� ������۟ɟ���#� 5��Y�G�}�k����� ůׯ������1�� U�C�y�g�������ӿ ������	�?�-�O� Q�cϙχϽϫ����� ����;�)�_�M߃� ��?��߿�i������ %��I�7�m�[�}�� �����������!���E�/�  e�i�� i�}�i��$T�BJOP_GRP� 21��  ?�i�i	������9�� � Y���� �����y���i� @e����	 �CB  ��C����5G�U	i�C 2BH  A�/���D�,��bB�* q�$�7C�� ���c�ad��i�A �EG+��a	���D/�D<Ky/�/ /#/�/�/��	? ?�/�/T?f?%?o?a	 �?�?�?�?�?�?�?O )OO!OOO�O[OO�O@�O�O�O�O_g�i��1Q�E	V3.�00��md45��*[P��d�i_tW� G/� G�7� G?h G�G8 GO G�d� Gz  G��� G�| G��: G�� G��� G�t G��2 G�� G�ݮ G�l G��* G�� H�S�RF� F�@ F+� F�K  Fj` F� F�Q � �GX �R�Q^�� Gv G����S�4 G�� �G�� G�\ �G� =L��/=#�
]Ae�JQs�Yokbi�oo��o��ESTPARb�P]����HR�`ABLE 1	���C`i��h�g ��di�g�hn i�h�Tp�g	�h
�h�hT�ei��h�h�h�Da�cRDI�o����o!3EWu�tO ��{����+��b	S��� �z���� "�4�F�X�j�|����� ��ğ֟�����0� B���Āȏ���g��l� ~�����N`r����x�bi�NUM  �1���	 �q� C`D`�b_CF�G 
R���@���IMEBF_T�T�a�����`��VE�RBc������R {1�k 8f_�i�d�� P���  ���%�7�I�[� m�ϑϣϵ������� ���!�3�|�W�i߲�@�ߟߵ�������A�����MD3�E���� k�}��V_I8����INT����b��T1�#�5� B��8O�a���_TC�����$�P����9�RQH��Դ_L���@˵��`MI_CHA�N�� ˵ nDB/GLVL��˵�a�q ETHERADW ?�e� ��`������hq R�OUT��!P�!�#ASNMA�SK�˳�255.GS}��GS��`OOLOFS_�DI�P�%�	OR�QCTRL ޻7��o-T/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?s<�/�?�?�?�cPE_�DETAI��P�GL_CONFI�G R�b����/cell/$�CID$/grp1�?4OFOXOjO|O2��
�O�O�O�O�O_ �O%_7_I_[_m___ �_�_�_�_�_�_�_�_ 3oEoWoio{o�oo�o �o�o�o�o�o/A Sew�*�� ������}�O� a�s���������?я������*�<�N� `����������̟ޟ m���&�8�J�\�n� ��������ȯگ�{� �"�4�F�X�j����� ����Ŀֿ������ 0�B�T�f�x�ϜϮ� �������υ��,�>� P�b�t߆�ߪ߼��� ������(�:�L�^� p������������ ��@�Us�er View �"I}}1234567890C�U�g��y�������. C����)�26���+@=Oa����0�3�� �����	h*��4�cu�������5R/)/�;/M/_/q/��/��6 /�/�/�/??%?�/F?��7�/?�?�?�? �?�?8?�?��8n?3O EOWOiO{O�O�?�O�B� lCamera4�*O�O_ _)_;_M_+�E�Ow_ �_�^A��_�_�_�_�_o)  �F���O_o qo�o�o�o�o`_�o�o Lo%7I[m�O��F�	��� ��%��oI�[�m�� ������Ǐُ돒�w Q��7�I�[�m���� 8���ǟٟ$����!� 3�E�W����w+k🥯 ��ɯۯ�����#�5� G���k�}�������ſ l��E�)Z��!�3�E� W�i���ϟϱ����� ������/�ֿ�wm9 ��{ߍߟ߱�����|� ����h�A�S�e�w� ���Bߤw!I2����� ��/�A���e�w��� ���������������9��HZl~� �I������� @2DVhz	J	�E0 �����/ �3/E/W/�{/�/�/ �/�/�/|��@�Ky/ .?@?R?d?v?�?//�? �?�??�?OO*O<O NO�/�EBk�?�O�O�O �O�O�O�?_*_<_�O `_r_�_�_�_�_aO� �{Q_oo*o<oNo`o _�o�o�o�_�o�o�o &�_�U��or �����so�� �_8�J�\�n����� 9�U��)�ޏ���� &�8��\�n���ˏ�� ��ȟڟ������U� ��J�\�n�������K� ȯگ�7��"�4�F�xX�j��  � ������Ͽ�����)�;�M�_�    o�w��ϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w������������c�  
�( � 荰( 	 ��;)_M �q�������%��� � ��j|����� ��/�Y6/H/Z/ �~/�/�/�/�/�// �/? ?g/D?V?h?z? �?�?�/�?�?�?-?
O O.O@OROdO�?�?�O �O�OO�O�O__*_ <_�O`_r_�_�O�_�_ �_�_�_oI_&o8oJo �_no�o�o�o�o�oo !o�o"ioFXj |���o���/ ��0�B�T�f���� �����ҏ����� ,�s���b�t���͏�� ��Ο����K�(�:� L���p���������ʯ �� ��Y�6�H�Z� l�~���ׯ�ƿؿ� 1�� �2�D�V�hϯ� �Ϟϰ���������
� �.�u�R�d�v߽Ϛ߀�߾�������;�@� �#�5�G���� ��0frh�:\tpgl\r�obots\am�100id\arc_mate_���_1450.xml�����������`�0�B�T�E���Y� ~���������������  2D[�Uz� ������
 .@WQv��� ����//*/</ SM/r/�/�/�/�/�/ �/�/??&?8?O/I? n?�?�?�?�?�?�?�? �?O"O4OK?EOjO|O �O�O�O�O�O�O�O_ _0_GOA_f_x_�_�_ �_�_�_�_�_oo,ot>n`��� �k�<< i�?�>k�o>oyo�o�o �o�o�o�o�o5- O}c���������1�?��$T�PGL_OUTP�UT I�I�/ a`i�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��i��a`�6�2345678901A�S�e� w�������?�>�ʯܯ � ��$���(�Z�l�~�����:�}��Կ� ��
�ϴ�ƿR�d�v� �ϚϬ�DϺ������ �*���8�`�r߄ߖ� ��@�R�������&� 8���F�n����� N��������"�4��� ��j�|���������\� ����0B��P x����Xj� ,>P�^� ����f�// (/:/L/�A�}\a�/@�/�/�/�/�/�-@co�?#?ij ( 	 &�X?F?|?j?�? �?�?�?�?�?�?OO BO0OfOTO�OxO�O�O �O�O�O_�O,__<_@>_P_�_t_�_4��_` xf�_�_�]�_o*oo No`o.��_�o�o=o�o �o�o�o!o%W �oC��y��3 ����A�S�-�w� ���q���яk���� ��=�����s���� ����������a�'� 9�ӟ%�o�I�[����� �����ٯ#�5�� Y�k�ɯS�����M�׿ �ÿ��}��U�g� ϋϝ�wω���1�C� 	�ߵ�'�Q�+�=߇� ���ϝ���i߻��� ��;�M��5���o� ��������_���7� I���m��Y������ %�������3 i{����K�����/�R�$T�POFF_LIM� �P��Qy��JN_SVN�  �$`P_�MON �U)b��2�%J�STRTCHK ��U`/hVTCOMPATu��dVWVAR ��"(y �� :/Y��J_DEFPRO�G %�%�MAInOLDA�DURAQ/�_D?ISPLAYU��j"INST_MSwK  �, �*?INUSER��$�LCK�,�+QUI�CKMEN"?�$S7CREA0�U "?tpsc�$�!�\0a9`r0_v9ST��`RACE_C_FG �"$uY	C$
?��8?HNL 2y*�P�1)+ O"O'O9OKO�]OoO�O�O�J�5IT�EM 2K ��%$12345�67890�O�E � =<�O_*_2S G !8_@[L �O �_C#�O�_
_�_�_@_ �_d_v_?o�_Zo�_jo �oooo*oDoNo�o roDV�oz�o�o |&��
�n� ���:�������� "�ʏF�X�!�|�<��� `�r�֏����L�՟0� �T� �&�8���D��� ҟ�^����گ�P� �t������4�ί�� �����(�:��^�� ��B�Tϸ�j�ܿ� ���6���ߎ�~ϐ� �ϼ���@��ϖ߼��� 2���V�h�z��ߞ�J� p���ߎ�
��.��  �d�$�6���B����� ����������N�  r���M��h��x� ��8J\�� ,Rd���� ��F//|$/� �{/��/��/�/0/��/T/f//?�4S�2|�?4:�  �B�4: �1�?�)
 ��?�?�?�?c:UoD1:\�<��F1�R_GRP 1��K� 	 @� :OLK6OlOZO�O~O�O�N��@�O�J�A��?_�O7_"U?�  R_d[N_�_r_�_�_ �_�_�_�_�_&ooJo�8ono\o�o�o�o�o	�5�o�oD3SCBw 2P; =_ :L^p������:<UTORIAL P;�?�?7�V_CONFIG  P=�1�?�?t��$�OUTPUT �!P9e��� ��ď֏�����0� B�T�f�x�����b��� ğ֟�����0�B� T�f�x���������ү �����,�>�P�b� t���������ο�� ��(�:�L�^�pς� �ϦϷ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r �������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ N�`����/??&?8? J?\?n?�?�?�?�?�? ��?�?O"O4OFOXO jO|O�O�O�O�O�?�O �O__0_B_T_f_x_ �_�_�_�_�_�O�_o o,o>oPoboto�o�o �o�o�o�_�o( :L^p���� ��o� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶���|�Ͻ(����� �����6��/Z�l�~� �ߢߴ����������  �2��V�h�z��� ����������
��.� @�Q�d�v��������� ������*<M� `r������ �&8I\n �������� /"/4/F/Wj/|/�/ �/�/�/�/�/�/?? 0?B?S/f?x?�?�?�? �?�?�?�?OO,O>O O?bOtO�O�O�O�O�O �O�O__(_:_L_]O p_�_�_�_�_�_�_�_  oo$o6oHoY_lo~o �o�o�o�o�o�o�o� 2DS{�$TX�_SCREEN �1"����}�S�������Bք1� C�U�g�y������� ӏ���	����?��� c�u���������4�� X���)�;�M�_�֟ 蟕�����˯ݯ�f� ���7�I�[�m���� ���,�ٿ����!� 3Ϫ���i�{ύϟϱ� ��:���^���/�A��S�e��ω��$UA�LRM_MSG k?sy��p �� Vj��������"��F� 9�K�i�o����������SEV  �����ECFoG $su}q�  Ve@�  }AJ�   B�Vd
 ��]csu}��� �������������1?&�GRP 2�%0� 0Vf	 �g����I_BB�L_NOTE �&0�T��#l]bxp_a<�?DEFPRO��Z�� (%��_` �*N9r]� ������/��FKEYDATA� 1'sys p 	?�Vfvy/�/b/�/�/�*,(�/�/Vd�([ INST� ]�/�.  IR�ECTR�D?+?ND�=2T?V? CHOI�CE?�?[ED�CMD�?�?� ORE0FO�?�?O*O ONO5OrO�OkO�O�O��O�O�O_�O&_8_� ��/frh�/gui/whi�tehome.png9_w_�_�_�_�_{�PVinstb_��_oo(o:o�W  >QUdirec�U�_�o�o�o�o�oVhin aj�o);�oXfchoicaS�o�������PPVedcmdo��'��9�K��VPVarwrg�o��������Ϗ Vx����"�4�F�X� �|�������ğ֟e� ����0�B�T��x� ��������ү�s�� �,�>�P�b�񯆿�� ����ο�o���(� :�L�^�p�GUuϜϮ� �����������,�>� P�b�t�ߘߪ߼��� ���߁��(�:�L�^� p�����������  ���$�6�H�Z�l�~� ������������� ��2DVhz� �����
� @Rdv��)� ���//�</N/ `/r/�/�/%/�/�/�/ �/??&?�/J?\?n?Ѐ?�?�??[�;�>JP����?�? �=�? O2OF,_cO _�OnO�O�O�O�O�O __�O;_"___q_X_ �_|_�_�_�_�_�_o �_7oIo0omoTo�o�o ���o�o�o�o!0? EWi{���@ �����/��S� e�w�������<�я� ����+�=�̏a�s� ��������J�ߟ�� �'�9�ȟ]�o����� ����ɯX�����#� 5�G�֯k�}������� ſT������1�C� U��yϋϝϯ����� b���	��-�?�Q��� u߇ߙ߽߫����߸o ��)�;�M�_�f߃� ����������~�� %�7�I�[�m������ ��������z�!3 EWi{
��� ����/AS ew����� �/�+/=/O/a/s/ �//�/�/�/�/�/? �/'?9?K?]?o?�?�? "?�?�?�?�?�?O�? 5OGOYOkO}O�OO�O��O�O�O�O__���![������J_\_n]F_�_�_|V,�o�_�o�_�_o-o oQo8ouo�ono�o�o �o�o�o�o);" _F�j���� �����7�I�[�m� ����O��Ǐُ��� �!���E�W�i�{��� ��.�ß՟����� ��A�S�e�w������� <�ѯ�����+��� O�a�s�������8�Ϳ ߿���'�9�ȿ]� oρϓϥϷ�F����� ���#�5���Y�k�}� �ߡ߳���T������ �1�C���g�y��� ����P�����	��-� ?�Q�(�u��������� ������);M _�������� l%7I[� ������z /!/3/E/W/i/��/ �/�/�/�/�/v/?? /?A?S?e?w??�?�? �?�?�?�?�?O+O=O OOaOsOO�O�O�O�O �O�O_�O'_9_K_]_ o_�__�_�_�_�_�_ �_�_#o5oGoYoko}o��of��k�f�����o�o�m�o �f,�C�g N������� ���?�Q�8�u�\� ������Ϗ���ڏ� )��M�4�q���b��� ��˟ݟ��o%�7� I�[�m���� ���ǯ ٯ������3�E�W� i�{������ÿտ� ���Ϭ�A�S�e�w� �ϛ�*Ͽ�������� ߨ�=�O�a�s߅ߗ� ��8���������'� ��K�]�o����4� ���������#�5��� Y�k�}�������B��� ����1��Ug y�������� 	-?Fcu� ����^�// )/;/M/�q/�/�/�/ �/�/Z/�/??%?7? I?[?�/?�?�?�?�? �?h?�?O!O3OEOWO �?{O�O�O�O�O�O�O vO__/_A_S_e_�O �_�_�_�_�_�_r_o o+o=oOoaosoo�o �o�o�o�o�o�o' 9K]o�o��������� �}�� ���*�@<�N�&�p���\�,n� ��f�׏������1� �U�g�N���r����� ���̟	���?�&� c�J������������ ���)�;�M�_�q� �������˿ݿ�� ��%�7�I�[�m��� �ϵ��������ό�!� 3�E�W�i�{ߍ�߱� ����������/�A� S�e�w������� ��������=�O�a� s�����&��������� ��9K]o� ��4���� #�GYk}�� 0����//1/ �U/g/y/�/�/�/� �/�/�/	??-???�/ c?u?�?�?�?�?L?�? �?OO)O;O�?_OqO �O�O�O�O�OZO�O_ _%_7_I_�Om__�_ �_�_�_V_�_�_o!o 3oEoWo�_{o�o�o�o �o�odo�o/A S�ow����� �r��+�=�O�a� ���������͏ߏn� ��'�9�K�]�o�F �q��F ��������������̖,ޯ#�֯G�.�k� }�d�����ůׯ���� ��1��U�<�y��� r�����ӿ����	�� -��Q�c�B/�ϙϫ� ����������)�;� M�_�q� ߕߧ߹��� ����~��%�7�I�[� m��ߑ��������� ���!�3�E�W�i�{� 
��������������� /ASew� ������+ =Oas��� ���//�9/K/ ]/o/�/�/"/�/�/�/ �/�/?�/5?G?Y?k? }?�?�?x��?�?�?�? OO&?COUOgOyO�O �O�O>O�O�O�O	__ -_�OQ_c_u_�_�_�_ :_�_�_�_oo)o;o �__oqo�o�o�o�oHo �o�o%7�o[ m����V� ��!�3�E��i�{� ������ÏR����� �/�A�S��w����� ����џ`�����+� =�O�ޟs���������hͯ߯�0���0���
��.��P�b�<�,Nϓ�F� ����ۿ�Կ���5� G�.�k�RϏϡψ��� ����������C�*� g�y�`ߝ߄����߲? ��	��-�?�Q�`�u� ���������p�� �)�;�M�_������ ��������l�% 7I[m����� ���z!3E Wi������ ���///A/S/e/ w//�/�/�/�/�/�/ �/?+?=?O?a?s?�? ?�?�?�?�?�?O�? 'O9OKO]OoO�OO�O �O�O�O�O�O_��5_ G_Y_k_}_�_�O�_�_ �_�_�_oo�_CoUo goyo�o�o,o�o�o�o �o	�o?Qcu ���:���� �)��M�_�q����� ��6�ˏݏ���%� 7�Ə[�m�������� D�ٟ����!�3� W�i�{�������ïR� �����/�A�Яe� w���������N����@��+�=�O�&PQ���&P����zόϞ�v����Ϭ�, ��߶�'��K�]�D� ��hߥ߷ߞ������� ���5��Y�k�R�� v������������ 1�C�"_g�y������� ��п����	-? Q��u����� ^�);M� q������l //%/7/I/[/�/ �/�/�/�/�/h/�/? !?3?E?W?i?�/�?�? �?�?�?�?v?OO/O AOSOeO�?�O�O�O�O �O�O�O�O_+_=_O_ a_s__�_�_�_�_�_ �_�_o'o9oKo]ooo �oX��o�o�o�o�o�o o#5GYk}� ������� 1�C�U�g�y������ ��ӏ���	����?� Q�c�u�����(���ϟ ������;�M�_� q�������6�˯ݯ� ��%���I�[�m�� ����2�ǿٿ���� !�3�¿W�i�{ύϟ� ��@���������/� ��S�e�w߉ߛ߭߿�ږ`����`����������0�B��,.�s�&���~� ����������'�� K�2�o���h������� ��������#
GY @}d���o�� �1@�Ugy ����P��	/ /-/?/�c/u/�/�/ �/�/L/�/�/??)? ;?M?�/q?�?�?�?�? �?Z?�?OO%O7OIO �?mOO�O�O�O�O�O hO�O_!_3_E_W_�O {_�_�_�_�_�_d_�_ oo/oAoSoeo�_�o �o�o�o�o�oro +=Oa�o��� ������'�9� K�]�o�v������ɏ ۏ�����#�5�G�Y� k�}������şן� �����1�C�U�g�y� �������ӯ���	� ��-�?�Q�c�u���� ����Ͽ���Ϧ� ;�M�_�qσϕ�$Ϲ� �������ߢ�7�I� [�m�ߑߣ�2����� �����!��E�W�i� {���.������������/��$UI_�INUSER  ����P��  0��4�_MENHIS�T 1(P��  ( �]���(/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,153,1o�������)����631���ew�� �'-?7S��
��.�?edit���SOLDADORA,3!t����35GMAIN_XU_��/ /��,�GIR_HOME�x/�/�/����/�/�/�/??,? �/P?b?t?�?�?�?���D1��D?�?�?OO )O;O>?_OqO�O�O�O �OHO�O�O__%_7_ �O�Om__�_�_�_�_ V_�_�_o!o3oEo�_ io{o�o�o�o�oRodo �o/AS�ow ������?�?� �+�=�O�a�d���� ����͏ߏn���'� 9�K�]�o��������� ɟ۟�|��#�5�G� Y�k���������ůׯ ������1�C�U�g� y��������ӿ��� ��-�?�Q�c�uχ� ���Ͻ�������ߔ� )�;�M�_�q߃ߕ�$� �����������7� I�[�m��� ���� �������!���E�W� i�{�����.������� ����Sew �������� +��as�� ��J��//'/ 9/�]/o/�/�/�/�/ F/X/�/�/?#?5?G? �/k?}?�?�?�?�?T?��?�?OO1OCO.���$UI_PAN�EDATA 1*����yA�  	�} � frh/gui��Adev0.st�m ?_widt�h=0&_hei?ght=10�@�@�ice=TP&_�lines=15�&_column�s=4�@font�=24&_page=whole�@�UO1)  rim�O!_  �@8_J_\_ n_�_�_�O�_�_�_�_ �_o"o	oFo-ojo|o co�o�o�o�o�o�o1�� �  �   I}� 2_7I[m��o �(_����!�3� �W�i�P���t���Ï ���Ώ���A�(� e�w�^���y��{C �۟����#�5��� Y��}�������ůׯ >������1��U�g� N���r�����ӿ�̿ 	��-�?ϲ�ğuχ� �ϫϽ���"���f�� )�;�M�_�q߃��ϧ� ���߲������%�� I�[�B��f���� ��L�^��!�3�E�W� i������������� ����A(ew ^������� +O6s���� ������//h 9/��]/o/�/�/�/�/ /�/�/�/?�/5?G? .?k?R?�?v?�?�?�? �?�?OO��UOgO yO�O�O�OO�OF/�O 	__-_?_Q_c_�O�_ n_�_�_�_�_�_o�_ )o;o"o_oFo�o�o|o �o,O>O�o%7 I�om�O��� ���d!��E�W� >�{�b�������Տ�� ����/��S��o�o}�d�������ӟ���)����u�H�Z� l�~�����	�Ư��� ѯ� ��D�+�h�z� a�����¿Կ�����x��c�k�$UI_P�OSTYPE  ��e� �	 �[�*�QU�ICKMEN  �9�H�^�,�RE�STORE 1+��e  '�뿑r�����ϑrm �)�;�M�_� q�ߕߧ߹����߀� ��%�7�I���V�h� z��ߵ���������� !�3�E�W�i�{���� ������������ ��Sew��>� ����+=O as(��� �//'/9/�]/o/ �/�/�/H/�/�/�/�/ ?�?0?B?�/}?�? �?�?�?h?�?�?OO 1OCO�?gOyO�O�O�O�i�SCREy�?�~�u1sc���u2�D3�D4��D5�D6�D7�D8��A�CTAT5�� ����e"�USER��@�O�BT�@�CksT�C�T4�T5�T6�T�7�T8�Q*�NDO_CFG ,9�Xt�s�*�PD-QgY��None� *�^P_INF�O 1-�e`��0%�O,o�xo[o >oo�oto�o�o�o�o �o!EW:{�b��QOFFSET' 09�a�PC ��XO����/�&� 8�e�\�n��r����� ȏ�����+�"�4�F� ���ϒ�����
��ڟ��xUFRAME � PD�V�QRTOL_ABRT����s�ENB��G�RP 11�Ɋ�?Cz  A�u�s� �Qs���������ͯ߯���x�U?��Q.�MSK  B�a.�mN��%	i�%b����k�VCMR[�2�7�{#�R@	��Pfr1: S�C130EF2 Q*ݿ�PD�����T�&��5R@�Q?���@�p��ȇ� ɟ5�?�IH`�@rϟ�ı����8�屢A�RB���RB? B����RA #ի�Dߋ�h�7ߌ�w� �ߛ��߿���
�a��� @�+�=�v�)ߚ��ISIONTMOiU�B��U�����R8SﳸS�� j� F�R:\��\�PA\��� �� M�C�LOG�  � UD1�EX�5�RA' B@ ��x�I�r����I����PC �� n6  ��q�IFu�%��`���Z�  =����PD	 J�*�TR�AIN_���ǐ  dPp	�栲9�}(c��W� ������.�2@Rdv���_\�RE��:b�ʲ��/LEXE��;�{�Q�1-e��VMPHKAS/P�U�S����RTD_FIL�TER 2<�{ Ԓ��,�{/�/�/ �/�/�/�/�/??�� i/N?`?r?�?�?�?�?��?�?�?��SHIF�T�1=�{
 <��q�JODU)OOO�O _OqO�O�O�O�O�O�O _<__%_r_I_[_�_�_	LIVE/�SNAPesvs�fliv.�_���� �pU�P�Rmenu�_�_�_Woio�@b	E��>IO�EM�O��?�� ��$�WAITDINE#ND��+��dO?�"���g���oS�iTI]M@���<|G�o ^}�o�{az/azN�hRELE%!@��dx�����a_ACT�Pp�K�E�� @d��ko���E�RDIS��PA��`V_AXS-R�p2Ab������Vp_IR  �j 	��)�;�M� _�q���������˟ݟ ���%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ�����n��XVR�aB���$ZABCp1�C� ,N f�2�ϵ�ZIP��D��e������ύ�M�PCF_G 1E�ٍ0J��=��S�F8ىX�`# �c��n��<90 ��`��S�|��ߠ�?�}� �����S��$�z�8�x���� ��� ��������
�4�M����G��JÛ�YLI�NDK!Hً ���� ,(  * ��������������� ��);M��p ���{���  U6��lS��w�����Y�2Iه]� �)�#/3, ���\/G/�/��/�/ڄ��!A�c�SPHERE 2Ju��*?z�/<?#?`? ��/�?�?$�?k?Q? O�?&OO?\OnO�? �?�OO�O�O�O�OEO�"_4_F_M�ZZ/� ǘf