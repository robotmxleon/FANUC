��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����DRYRUN_�T  4 �$'ENB  �$NUM_POkRTA ESU@�$STATE }P TCOL_���PMPMCmGR�P_MASKZE�� OTIONNLOG_INFON�iAVcFLTR�_EMPTYd ?$PROD__ L ��ESTOP_D�SBLAPOW_�RECOVAOP�R�SAW_� G� %$INI�T	RESUME�_TYPENDIST_DIFFA $ORN41� 8d =R��&J�_  4 u$(F3IDX�̈_ICIfMI/X_BG-y
�_NAMc MO�Dc_USd�I�FY_TI� �MKR- � $LINc  � "_SIZ�c�� �. X� $USE_FLC 3!�:&iF*SIMA7#QC#Q�Bn'SCAN�A�X�+IN�*I��_oCOUNrRO( ���!_TMR_V1A�g#h> �ia �'` �����1�+WAR��$�H�!�#N3CH�PE�$O�!�PR�'Ioq6�$�$CLASS  �����1��5z��5�0VERS���7  {�ץ1IRTU� ��?�0'/ �5+5��������0BF�0�1E��%�1 9O��5OnO�����5vI2�; vO �O�O�O__%_7_I_ [_m__�_�_�_�_�_��O)W?�8�0 ��j�0*o<orNi�� � 2�9?  4%�_�o��AA�o�o�o�o��o%7[��@ �AM�=�������dcs�yjc$"P+ uk"K�0��U�A`�XA�1�0$N ��������Џ��� �*�<�N�`���FA u�A������ʟܟ�  ��$�6�H�Z�l�~�̘4L!�C� 2ulu�ۯ��� �#�5�G�Y�k�}��� ����t�ͯ���
�� .�@�R�d�vψϚϬ� ��ɿ������*�<� N�`�r߄ߖߨߺ��� ������&�8�J�\� n����������� ���"�4�F�X�j�|� �������������� 0BTfx�� ������, >Pbt���� ����/(/:/L/ ^/p/�/�/�/�/�/�/ �/rv