��   v1�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����UI_CONF�IG_T  � E$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]5�ODE�
6CWFOCA �7C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"�%�!BA�!j ��!�BG�#�!hINS�R$IO}7P}M�X_PKT?$IHELP� {ME�#BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�<ST]Yf2$Iv!_Gv!k FKE�E ��8C &USTO}M0 t @;AR$@PIDDbB�ChD*PAG� ?�^DEVICEބISCREuEF���}GN�@$FwLAG�@3&��1  h 	$�PWD_ACCES� =EFB�S�:1�%)$LABE�� $Tz jp�@�32R�	c&�USRVI 1  < `'R*'R��(QPRI�mx� t1�PTRIP�"m�$$CLA�@? ����Q��eR��R�P\ SI���W  ;�׸QIRTs1�_��P'2 L17�L�1A�R�	 ,���?���a�P$bda��>a���`�  �����
 ��'/�SOFTPb@/G�EN�1?CURR�ENT=>�A,18,1lo�o�o�o�o� �o�o,95,2��o?Qcu �(5�`w�����)q9�G�Y� k�}����s�oˏݏ�������E,381�oN�`�r�����Q ������ӟ���	��� -�?�Q�c�u������ ��ϯ�����)�;��M�_�q�����a_TPTX��&����˿` s�����$/softp�art/genl�ink?help�=/md/tpm?enu.dg��2� D�V�h�!��Ϟϰ��� ����u�
��.�@�R� d���uߚ߬߾����� �߃��*�<�N�`�r�V����Q[fAfc��($��������������Qa:� <cI�<c:�8����zc��\a?d�����  ��	���K�����`�[`^�W`  ��� ���SQB 1��XR \���_�� ;REG VED��F�Xwholem�od.html	s�ingl}do�ub�tri�p�brows�t�Y�� CUgy��C-|gydev.s��l/� 1,	t 0/�/��/�/�/�m/�/�/�/�/?8?� �PP?b?t?�?�?��?�?�?�?�?�6 @ L?!O3OOWOiO{OJF ;	3?-?�O�O�O�O�O 	__-_?_Q_c_u_�_ �_�_�_�_�_�_�o o3oEoWoio{o�o�o �o�o�o�o�o/ ASewE?��� ����0�B�T�OO x���Y�k���ҏ�O�O ���'�9�b�]�o� ��������ɟ���� �:�5�G�og�a��� ����ůׯ����� 1�C�U�g�y������� ��ӿ�� �2�D�V� h�zόϞϰϫ����� �����.����ݿv� q߃ߕ߾߹������ ��%�N�I�[�m�� ���q��������� !�3�E�W�i�{����� ����������/ ��j|����� ���0B# x�A�S�9��� �//'/9/b/]/o/ �/�/�/�/�/�/�/�/ ��??G?Y?k?}?�? �?�?�?�?�?�?OO 1OCOUOgOyO�OY�O �O�O�O_ _2_D_V_ h_c�_�_m__�_�_��Z�$UI_TO�PMENU 1��PaR� 
da�A)�*default��O�M*lev�el0 *�K	 #Ho60�o/o�o��btpio[23�]-8tpst[1�h�o�o�oko}o(=�h58E01_�l.png</6menu5^yUp�qC13^zr]z}t4�{l)q����
�� .�@�R��B�{������ÏՏd�pri�m=�qpage,?1422,1܏� '�9�K�]�h�������з�ɟ۟j���class,5��+��=�O�a�l���13�h�����¯ԯ�m���53�"�4�F�X�j�m���8����� ɿۿ�l��#�5�G�Y�kϖI`a.o�πRm��+q������ft�y�m�o�amf[0��o��	�c[164�gf�59�h+q�ߣ�yx2��}�ҙz ��w]{��s����n� ������������ �"�4���X�j�|�������A���2���� /A���w�� ��N`�� $6H��	�1\��Ъ��M���ainedi��//)/�;/M/H�conf�ig=singl�e&��wintp ��X/�/�/�/�/�Ja ���/?Se?%��E? W?i?|?�?�?�?�?1? �?�?OO/OAOSOeO wO��O�O�O�O�O_ _M�>_P_b_t_�_�_ '_�_�_�_�_oo�_ (oLo^opo�o�o�o5o �o�o�o $�oH Zl~��1�� ��� �2��V�h� z�������?�ԏ���
��.��N��d���@�����ϑO��5�s�̟�'�ٗuݤ���  �����3��ڂ�����̩6ٯu7�F�X� 1�C�U�g�y�ď���� ��ӿ������-�?ϠQ�c�uχ�f"\1 k��������	��-� ?�Q�c�u߇�߽߫� ��������Z�M�@_�q���$�6�6����������d$�74$�U�g�y������,�C���5	TPTX�[2096��4��2�46�������18@"4F��0��25��1��i���tAvԡ����0��1���C:l$treeviewy#��3C�&dual�=o�81,26,4$�����/ ///A/S/e/��/�/ �/�/�/�/&�;x�53��E�O?a?s? ~/�?�?�?�?�?�?�? O'O9OKO]OoO�/?:�1%?�2���O�O��O �6�O.�edit��O�OT_f_x_ '�w5�1_CS�_�_�_ o��o4o�<o�Uo !{o�o�o�o�o�o�o go/ASew �������� "�4�F�Oj�|����� ��ďS������0� B�яT�x��������� ҟa�����,�>�P� ߟt���������ί]� ���(�:�L�^�� ��������ʿܿk� � �$�6�H�Z�	oo�� ?o����������  �1�C�U���aߋߝ� ����������	��@� R�d�v�������� ������*���N�`� r�������7������� &8��\n� ���E��� "4�Xj|�� ��S��//0/ B/�f/x/�/�/�/�/ oρ��/��?���=? O?a?s?�?�?�?�?)? �?�?OO(O9OKO]O oO1�O�O�O�O�O _ _]/6_H_Z_l_~_�_ _�_�_�_�_�_o�_ 2oDoVohozo�o�o-o �o�o�o�o
�o@ Rdv��)�� ����*��N�`� r�������7�̏ޏ�� ��&��/�/\�?�� �?�O����ǟٟ��� �!���-�W�i�{��� ����ïկ�O��0� B�T�f���x������� ҿ������,�>�P� b�t�ϘϪϼ����� �ρ��(�:�L�^�p� ��ߦ߸������� � ��$�6�H�Z�l�~�� �������������� 2�D�V�h�z���:�H��*defaul�t��j�*level8�M��	��� tpst�[1]	KyPtpio[23R6HuP�����menu7_l�.png��1	3�	5
��41u6�
�w� ������// +/=/O/�s/�/�/�/�/�/�/n"pri�m=�page,74,1�/?-???�Q?c?n"�&class,13h?�?�? �?�?�?u?�25�?"O 4OFOXOjOm#|<O��O�O�O�O�O�/218?)_;_M___q_|O�26x_�_�_�_�_�_���$UI_US�ERVIEW 1�J�J�R� 
�ED�IT,Weld �DATA s�d_oublej���_~�medit1@eo�o�o�o�okj�&95P�o,> �o�ot���p�0c�STATUS,P{OS@ftripMo _oqo�,�>�P�b��Yy2m�����ÏՏx�33_��1�C� �P�y�t������˟ ݟ����%�7�I�[� m��������ǯٯ�� ���
�|�E�W�i�{� ��0���ÿտ���� ��/�A�S�e�w�"��� �Ϩ��������+� ��O�a�s߅ߗ�:߻� �������ϸ�"�4� ��X�������l� �����#�5���Y�k� }�����L������D� 1CU��y� ����v�	 -?��L^p�� �����/)/;/ M/_//�/�/�/�/�/ v�/�/�/n/ ?I?[? m??�?4?�?�?�?�? �?�?!O3OEOWOiO? vO�O�OO�O�O�O_ _�OA_S_e_w_�_�_ >_�_�_�_�_o�R