��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A   �����
�WVAMP_�T   �$X1  $kX2AY@ /�FC5  �$2ENBA $�DT  / _�R2 d EN�ABLEDnSC�HD_NUMA ���/ CFG5�� $GRO�UP�$z ACC�EL@�G$MAX_FREQ�z2 L�DWEL��DEBUG�PRwEWSOUT�>PULSEA�SHIFt 7TY�P4$USE_�AEF} 4$G{DO�  f0 r?�Np�WEAVE_TS�K �V�_G�P�SUPPOR�T_CFnCNV�T_DONE �p }k}GRP G2r�� _� ��$� TIME�1�o$2'EX�T� (1#&(MODoE_SW�CO3 �SWIT � �P�HAX6  4 m� ECC$��TERMNnP�EAKno!AL ? \ � �!�I�$�!N_=VSTAR�#!�r"��"�%�C�YCL42 
� $/ � Tv"�b $CUR_R�EL_� �!��/ W�PR5 � 
�$CEN� _RI�3RADIU��XIz ] Z�IMUTi!$E�LEVATION�g5� N�CONTINUOe2q �MoEXAC=PE�8��6  H~ ��UENCYA�I�TUD4�2RIG�HC�2LEBL_�ANG1 �O�TF_� 	��  $3A�bE�T��n3C!�$ORGjHFB)KjH��P��C�.�DLDW�HR�E�_�3�B�C��D�B�Cp�@�D�A�CCHG�G�	Q�F	Q�F	Q�FINC�G=Q�F=Q�F=Q�F؃AVCPYC� _T��\#�Y~P#�@SY��H)@�UPD�"0n�$$CL�ASS  �����Q��8 �P�PV�ERS�1�W�  ���QIRTUAL�_�Q0� 2�X� � ��?��@�  HaDae�TWoio�{o�o�o`)dN 2� 3k Hf��=uHe@O�Hi�o�Nc)a� � e�� E`��`9t
��2�  �����=������4s �����jpYq��w�r��Dq��xat��ujp `��i.�5t8q�q�2�b�t���
�9x��������̏�ҏ���Sb)a�  2�3k
TDacSI�8� �����j0h�?m�'�� ��l�D�����Ca��l� ���k��� �2�D�V��h�z��lFI�GURE 8�� o�v�Hal�f������ ��M�(�H��󈯎�࠿��Ŀֿ�T'CIR1��Pd� }�0�~�h�z�D�Z�l���0�v˜�~�����p ��$ߪjN�� Hp��4q�Ȓ���@ ��ʖD�M`g������ ����	��-�?�Q�c�u`�� �>q� �5)�ᐟ N`���ᬟ����˟�� ��M�_�q�������������kTriangle��z� h߾�M��Ɵ�ύ� �����/ L�&��g �n���	//-/ ?/Q/c/u/�}DVh z��/�/��9?K? ]?o?�?�?�?�?�?����� O�h��O2O DOVOhOzO�O�O�O�O �O�O�O
__.[�?._ O"O�_�_�_�_�_�_ �_oo&o8oJo\ono��mSCHEXTENB  =��ct�STATE 2�k |o�o�o ��gWPR �7�6�L}D�-�_OTOF 	8��@)0��q�q���v)��uA�ȫs�u@�  <#�
�?����mu�_GP 2w| ���d�v���� я㏡+