��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A   �����
�WVAMP_�T   �$X1  $kX2AY@f/�FC5  �$2ENBA $�DT  / _�R2 d EN�ABLEDnSC�HD_NUMA ���/ CFG5�� $GRO�UP�$z ACC�EL@�G$MAX_FREQ�z2 L�DWEL��DEBUG�PRwEWSOUT�>PULSEA�SHIFt 7TY�P4$USE_�AEF} 4$G{DO�  f0 r?�Np�WEAVE_TS�K �V�_G�P�SUPPOR�T_CFnCNV�T_DONE �p }k}GRP G2r�� _� ��$� TIME�1�o$2'EX�T� (1#&(MODoE_SW�CO3 �SWIT � �P�HAX6  4 m� ECC$��TERMNnP�EAKno!AL ? \ � �!�I�$�!N_=VSTAR�#!�r"��"�%�C�YCL42 
��� Tv"b �$CUR_RELq_� �!3WPR5� � 
$CE�N� _RI3RA�DIU�XI�z ] ZIMU�Ti!$ELEV�ATIONg5� N��CONTINU�Oe2q �MEXAC=PE�3�6 � H~ �UEN�CYA�ITUD<4�2RIGHC�2�LEBL_ANG�1 �OTF_�� 	�  1$3A�bET���n3C!$O;RGjHFBKjH���P��C��DLD%W�HR�E�_�3�B �C��D�B�C�@�D�A�CCHG�G	Q�F	Q8�F	Q�FINC�G=Q �F=Q�F=Q�F�AVCPYC� _T�\#�Y�~P#�@SY��H)@�UPD"0n��$$CLASS  ����Q���8 �P�PVERS��1�W  ����QIRTU�AL�_�Q0 2~�X�  ��{?��@�  Ha Dae�TWoio{o�o�o�`)dN 2 3k� Hf��uHe@O�Hi�oNc)a� � e� E`���H��$��
��2 � �����=�s����4s �����jpYq��w�r�� Dq��xat��ujp`���i.�5t8q�q�2�b�t���
�<q` �����@q����̏ҏ����Sb)a�  2�3k
TDaS1I�8� �����Cp5h�?m�'���� l�D�����Ca��l��� �k��� �2�D�V�h��z��lFIG_URE 8��o� v�Hal�f������� �M�(�H��󈯎����Ŀֿ�TCIR1��Pd�}��0�~�h�z�D�Z�l���0�v˜�~����� ߸�$ߪjN� @Hp��4q�Ȓ���@�� ʖD�M`g�������� ��	��-�?�Q�c�u���`�� �q� �5)�ᐟN` ���ᬟ����˟��� M�_�q�������������kTriangle��z�h� ��M��Ɵ�ύ�������/ L�&��g� n���	//-/?/ Q/c/u/�}DVhz ��/�/��9?K?]?�o?�?�?�?�?�?�� ��� O�h��O2ODO VOhOzO�O�O�O�O�O �O�O
__.[�?._O "O�_�_�_�_�_�_�_ oo&o8oJo\ono�m�SCHEXTEN�B  =��ctSTATE 2�k |o�o�o ~�gWPR 7��6�L}D�-�_OTF' 	8��@)0�q��q���v)��uA���s�u@�  <#��
�?����mu_�GP 2w| � ��d�v����я ㏡+