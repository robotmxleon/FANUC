��   F��A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A #  �����#�AMON_D�O_T   �$PORT_�TYPE  �@NUMJ/SG�NL7 L�$MIN_RAN}GI$MAXr�NOo ALxp V��~ �COUNT>J��AWE08 �� $AWn0ENBJ $�|G1LY_TIV�$WRN_ALM�STP�
�E��C�.�WT�C�
J�AFT_�CHGxAVRG�_INT��{SgAVE�YP1?ER_REG�Tw$WA� SIG�� OP��V/OLTS�����AMP�&AEx �#E_VL� �&D'>% I*f$� _�ANL�  �p 
$US0 S�_CMD � PRIORITY�"�UPPER� $�LOW�$�#$FgDBK�"�RAv ~�!SQ_AVG�#n�#SD_� CE� 8� ��$ �� � �LIN�!$ARC_ENABL�!|� 0DETEC�!~< ELD_SP�$?PD_UNI��!N92DIS�"�ID sIM�#�� l v1WFt2θ�CF�" � �$PS_MANU�F �2OD�EL�5PROCEySN0�0WFEEW0�ESC�2�2_FI�#1�1�1�7T _AOT�"�2I�6D�7DC`1�6L �"{2 � �CNV� 7   $EQ�zx�ODOU��2?@T�Bd  $~?C 2 kE�DD   , �� MM�!�$D� ��!2� $F� �B�4NuV7	JBSEL10�_NOJDATA�_s@�@ �2W�PpG
{M
�FWP�7 L@�L
 ��WIR_CLP4 L@AS�BU8  H $(4��R�4�YPREF� �U��_ECU��  �JB~ �S  � $BPEEPf#�}!SCH7 � �!��`�1e�#dPK*jFRE�Q.gULSwbSP�0fg2y�!hybl*g�F� AI6 �ZCoVG}�h p dD�e�e�`�	�a���dBVB�aZERqOy}uSLO]R�`NT�!P�cO	U\�93�L FORMA�0NAra�0J3	� D�cQWUX�WEIOEX7O4 �A�Wfx�ccpS_91IN�p� :1�U�p� FcAUG"t0LO�0�qP�!�G��R<�yADp;�STIC�@��pROBOT�A{DY�rERRO�SE��`S��p�!�TR��$S�CHD�OG_�@%��0_AOCTIV���I��C�01�2�q�O�TF7 � $
��P��x�nfpNCi0�c;� f0�*d;�*g0�7f;� 7i0�Fd;�Fg~�Td���TfUP�@�B�3PC�R7�� WS#TK��� =�Hr Ւ Ɓ%��00��2�X���0A~�3KIPTHE91�S;������PIKEf���0��0WWV�2t�E_�HO;0�0��PHKp-1���� RMT����SPTL�0p�3$Hz��SW��pd�$BBg1_ONL4�$B�2pf�bgF�WF�1e2_R`��zE"�!� _W;6~�AND1OFF��.�!ND2g�3g�R��S� �A� 9CEPM~� | $�0 �@g��e��*f��7b���Ff�TfADAP�T� G�CSENS��c��!ݒ��8 � 0?,2���"� �$�1b�!c�7cc�Fa |�Tac�^��'y��&l�T�&�!4�&5�&6�"p8�W�@�2 HOU�!��o � �SE �0�g4�Q�T<��6 �'��46�q56�0� %$CURR7�(��"HEATzP e@�!燰"j���i�p.��GAP�#Ti�XP�Y0��EHP��@��pDYS�@�!GP�0S�!�$���$GO� RI���AM�#/"�#�M��jAN3O�BE	FB ;�LHV1[5j�@�43;1 `H�V�PA�H�r���3��F1�� ��DPOSR 7� � 	� RSB �$��0G�m�b�O�J�X��O��DU�IW�"AXQl�2C,1L»"D����?3ܓRG�8  4�@P֋q]ִSGʦ�~�;A8�~8  $ $�@ �CL�$��s	-đ�>8 $ ;o2� ��"�ql��q��� 	PK�P��
��*���q��Ba��b�@4
�5�6:2K�3�0����FW�q�yB��ALAR�� �2��2�����:
�3�Q_R}���
�.44�F�+�PW,���_@ĸ�Ӕ] �������Qbwm��t���QDI�c�j���~pus�R�SIZ<���BOAR���1"]E7�]�\��h"0h"��ķ�$�VEND��I��DOEVIC��0D�Ӯ��MAJ��V�#I�N�(�$�uI"�vMA��pFI�0�BW���RE�� p �$��X�� ⡡��F&̀OR_R��C�^1�D4TO_��O5_Rf�pRS�Q'�OS�9��rUP� #N��S�0�`�=� �6���6��9PURGX��RKtSTFR�p&���A��.E�.E@�AED��P-��M%�BfMT�����eEM7� �Q�5���Z$�22�9���P駇��K�p�QAD9J�T��NEXT��r'_LE�c��P��X���M����aA��_�#IV���H�q�2�e#FL������P��U����0�8� ��TWTl[�CY�� �>�  �	`���`( �bTOTAL!_�Q�c���VI�p�WGWARo��U��A*��PY&1b�uKG@���'" A}�#N�p�  #1SCF�G�1�`LO!O�B:��P�Q�S!x@���GLOB�Pp�⣠� ��NOT�ы$0QI4�*��AVh�Y��$����������e��W_SHFJL�W�X�fkrI�0$�q �e�RY	���p�P��%�ʀLIMS`p�i�@�c7�UIF�e��APCOUPL>�R @ �p�ql��� �qUR�`uN��<�MMYm 0�u0�u�  �����USTOk�    x�0 �qp`� 
��SEMG�g��1! ,��MGX�Ag���NOzPR ���wa�"� ,/���Ȣ=6Ƞ��3T� )�RT���Y���0=����AHER� A�������'"݈{�� �����@���Q�L�� )BD ��2C���7B<�^i3_FIL@�W��7BUG_3SM ���ñF_F����Z�, �_4N SV@БTC�P��=Ҕ�DIO��������.a�TM�C��PA�Pq��q�w�x��q�_DYN�V�2Wԣ����KE�YV�GQׂ��F`��?�/B�{�_C��R�TOU���������CAL�Q0�`�� TIp1�P_y�R�T���@��A?2���$$CLASS  ������ ��� �-�S�B���  ����IRTUx�����AWAOY1��� 
��$�a
�K���n�2�f�[�[���g�
�?�������g��� ��������(�:��L�^�pςϑ�l�EXEu�`���������Ͽ �*�<�N�`�r߄ߖ�p�ߺߕ�r@S Rw���:����#�5�G� Y�k�}���������������l�NLG7 2x� �����E?��<1�6�`��e�� p`����{` 2�:�)��General Purpose��MIG (V�olts, 0)���� ����
AW�MGENL.VR�A*EGLM#G19��g�`�� ������'���������������C�NV 2	x��[����� 4aPzUh �����//� =/O/./s/�/\�/�/ b/�/�/�/?'??K? ]?<?�?�?r?�?��E �/�?O�?2ODO#OhO zOYO�O�O�O�O�O�O 
__�?@_R_�Ov_�_ g_�_�_�_�_�_�_o �_(oNo�?ro-_�o�o 3o�o�o�o�o8 J)nM_�{o� ����� �F�%� j�|�[�������֏� go���0�B�!�f�E� W���{���ҟ����� �,�>��b�t���� ����ί௿����� :�L�+�p����O��� ʿU�� �߿$�6�� Z�l�KϐϢρ����� ����ߵ�2�D�#�h� z�Yߞ�}ߏ��߳����
��NVWP 2�|	i\>�T 
���b�t���UST�OM 2|l  ��������h��	hd"���DEF�SCH R|��Q�<�b�@De�fault Schg���n��������� ��K"4� Xj��������
)�FBKLOG�1 @��T���  Ugy��12=O�����5LG_CNT � ����)�IOE�X 2�����A� ��C�]$@�������!�
Weld Spee%�~�IPM  d$ �/�/�/�/??(?:?~��OTF 2���A?�?�?�?�?�?�C8=�����@����?K)�PCR k2��pI�BH�?��BC!�FK<D7�������?�ffA�Z �A"��OFM"@�����/�O@O�"@�����WOELG��k%*_�F��0234567O8901JRUK%4_y_�_�_HIȩ_7]�O_OSRAM2��I�B�$�_oCRGS_EL R<�Q�� 	Proce�ss 1oSf2T�_oj3i�o4i��o5�-mlXS��R�o7��kn8i'l�"@��� �_);Es-B� �W�%�Volta+ge��qsfc%�Dw|!@]y��h��aWiore f�  s�$	� hc%[&t/�o DS�l*�<�N�`�r� ��������̏ޏ��� �&�]+zvd"�����  �#��E��Z"!��a��^/�� ��V���a�aɒ�Curren=t�Amp�=� ��l�eu���Q�c�u� ��������ϯ��� �)�;�M��W���a�� ���ឱ	q��)q��Iq ��R�͹ϧg�a�aA� �b-���-�	q-�)q-��VE!��\e�	q/?�����Z�%�� ����ϻ������PD�RuS R\zH�� jq��C�U�g����� gߩ߻�u߇ߙ��� ������]�o�)�;�M� ��������#��� ���k�}�7�I�[��� ��������1C�� I��Wi�� ����?Q /������/ /)/;/M+�U/g){/��/�/M/�/?cS2�S�^=R��b�S2UP�Yp^=�=�o�?�33H1>E0=OL��>I0h!�"�#�$�1t9�g��q�#?�v�#>��8�8CWIRE �2&M<�?�?h��>�3�>�G(�=�J*�ESCFG �G�A��Y���OOˎE7])COU�PL�0=k
0 �vkB`�D�^�L�[�O ZW�O�G_�OP_G_Y\>�HNB  ��Ec�&FUSTOM � =k
8ƙy�O&EE�MGOFF !�=kS��)BPCRg "�_�@���zqC{sUūMJo�\zt�f_oeo��
Cl�q� �1