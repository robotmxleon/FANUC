��   F��A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A #  �����#�AMON_D�O_T   �$PORT_�TYPE  �@NUMJ/SG�NL7 L�$MIN_RAN}GI$MAXr�NOo ALxp V��~ �COUNT>J �AWE08 �� $AWn0ENBJ $�|G1LY_TIV�$WRN_ALM�STP�
�E��C�.�WT�C�
J�AFT_�CHGxAVRG�_INT��{SgAVE�YP1?ER_REG�Tw$WA� SIG�� OP��V/OLTS�����AMP�&AEx �#E_VL� �&D'>% I*f$� _�ANL�  �p 
$US0 S�_CMD � PRIORITY�"�UPPER� $�LOW�$�#$FgDBK�"�RAv ~�!SQ_AVG�#n�#SD_� CE� 8� ��$ �� � �LIN�!$ARC_ENABL�!|� 0DETEC�!~< ELD_SP�$?PD_UNI��!N92DIS�"�ID sIM�#�� � v1WFt2��C�F�" � $�PS_MANUF� �2ODE�L�5PROCES�N0�0WFEEW0EsSC�2�2_FI#1p�1�1�7T _AO�"*�2I�6D�7DC1��6L �"{2 � C�NV� 7   $EQ�zxOD�OU� A<CT�Bd� $?C �2 �?@D�D   , �� MM�!$�D� ��!2 �$F� �B�4NV�7	JBSEL10_�NOJDATA_�s@�@ {"WP�pG
{M
�
�DW�P7 L@�L
� �WIR_C;LP4 L@A�SBU8  H Q$4��R�<4�YPREF� �U�;A_ECU��  �JB~ �S  / $BPEEPf#�}!SCH7 � �!��`�1�e#dPK*jFR;EQ.gULSwbSP�0fg2y�!h�yb*g�F�"AI6 �ZCoVG}�hp  dD�e�e�`�	�a��d�BVB�aZERO8y}uSLO]R�`NT�!P�cO	U\93|�L FORMA0�NAra�0J3	�� D�cQWUXW�EIOEX7'4 �A�WfxccmpS_91INp�� :1�U�p� FA1UG"t0LO�0�q�P�!�G��R<�A<Dp;�STIC�@�p�ROBOT�AD�Y�rERRO�S�E��`S��p�!T�R��$S�CHDO�G_�@%��0_AC�TIV���I�Cʯ01�2�q�OT�F7 � $ 
��P��x�nfpNCi0�c;�f 0�*d;�*g0�7f;�7i 0�Fd;�Fg~�Td��Tf�UP�@�B�sPCR�7�� WSTK��� =�Hr ՒƁ %��00��2�X���0�A~�3KIPTH�E91�S;������PIKEf���0�0�WWV�2t�E_HaO;0�0��PHK-18���� RMT����SPTL�0p�$�Hz��SW��pd�$BBg1_ONL4�$B�2pf�bgF�WF�1e2_R��0zE"�!� _W;6�A?ND1OFF���!�ND2g�3g�R�Sp� �A� �SEPM�? | $�0�@ g��e��*f��7b���Ff�TfADAPTz� G�CSENS��c��!ݒ��8 � 0?,2���"��$ �1b�!c�7cc�Fa|� Tac�^��'y��&l��&*�!4�&5�&6�"8��W�@�2 HOU�!h�o � �SE�0 �g4�Q�T<��6��'��46�q56�0� ?%$CURR7(�^�"HEATzPe@ �!燰"j���i�p��GAP�#Ti�XPY0���EHP��@��pDS��@�!GP�0S�!�$���$GO� RI����AM�#/"�#M䩰jAN3O�BEFB ;�LHV1[5j�� 43;1 `H�V�PA�H�r���3��F1�� [@�/�SR 7 �+ 	� RSB�$�� 0G�m�b�O�J���O��DU�IW�A�XQl�2C,1L�"D�����?3���8 � 4�@P֋q]ִSG�ʦ�~�;A8�8  $ $�@�CL�$ć�s	۔��8 $ ;o2� �"�ql�0�q��� 	PK�P�� 
��*���q�BPa��b�@4�5�6:2K�3���&��FW�q�B��ALAR���2��2@�����
�3�Q_R}��
�.4�4�F�+�PW,���_ @ĸ�Ӕ]���� ���Qbwm��t���QDI�c�j��~pus��R�SIZ���BGOAR���1]E7�]�\�h"0h"��ķ�$VEN�D��I��DEVI�C��0D����MA5J��V�#IN�(�$�uI"�vMA��p�FI�0�BW����� p $��X��h ⡡��F̀OR_R���C�^1D4TO_l��O5_R�pRS<�f'�OS�9��UP� #N�:��0 �`�=� �6��6��9�PURG��RKtS�TFR�p&���A ��.E�.E�AED��P$-��M%�fMT�����eEM7��Q�5��� Z$�22�9�P駇��K��p�QADJ�T��NsEXT��r_LE�c"��P��X��M����aA��_�#IV���1H�q�2�eFL������P��:����0�8� ̀�;�WT[�CY���  �aE�  �	`��`( ~�bTOTAL_�Qȑc���VI�p�WWARo��U��A*�P1Y&1b�uKG����'" A}�#N�p { �SCFG�1wz�LOO�B:��P�Q�S!@���GLOB�P�⣠ܽ ��NOT��$b0QI4�*��AVh�Y��$��������e���W_SHFL�W�X�fkrI�$�q �e�RY	��оP��%�ʀLIMS`�i�@��c7�UIF�e�A�PCOUPL�R @ �p�q���[ �qUR�`N��<�MMYm �u0̼u�  ����US�TOk�   � x�0 �qp` 9
$�waEMGg��17! ,��MG�Ag���NOzPR ����|wa�"� ,/� ��Ȣ=6Ƞ��3T� )�RT���p�=����AHER�A��� ����'"݈{������ �@���Q�L��)BD���2C���7B<�i3_�FIL@�W��BU�G_3SM ���ñF�_F����q�, _4N& SV@БTC�P��8=Ҕ�DIO����`���.a�TM�C��PA�Pq��qw�x�<�q�_DYNV�2qWԣ����KEYV�!GQׂ��F��?�X/B�{�_C��R�TOU�����Б���CAL�Q0�`� ThIp1�P_y�RT����@��A?2E�$�$CLASS  _����� ��&� �-�SB����  �=��IRTU�����AWAOY1��[�$�
�K����n�2�f�`[�[���g�
�?��� ����g��������� ��(�:�L�^�pς���l�EXEu�`��� ������Ͽ�*�<�N� `�r߄ߖߨߺߕ�r@S Rw���:��� �#�5�G�Y�k�}����������������~l�NLG 2x�S �����?��<1�$6�`��e��� p`�����{` 2:��)�Gene�ral Purp�ose�MI�G (VoltsK, 0)��� �����
AWMGEN�L.VRA*?EGLMG19��g�`��������'� ��������������CNV 2�	x��[������ 4a PzUh���� �//�=/O/./s/ �/\�/�/b/�/�/�/ ?'??K?]?<?�?�? r?�?��E�/�?O�? 2ODO#OhOzOYO�O�O �O�O�O�O
__�?@_ R_�Ov_�_g_�_�_�_ �_�_�_o�_(oNo�? ro-_�o�o3o�o�o�o �o8J)nM _�{o����� � �F�%�j�|�[��� ����֏�go���0� B�!�f�E�W���{��� ҟ������,�>�� b�t��������ί� ������:�L�+�p� ���O���ʿU�� � ߿$�6��Z�l�Kϐ� �ρ����ϯ���ߵ� 2�D�#�h�z�Yߞ�}�����߳���
��NV�WP 2|	i\>�T 
��b�t�����USTOM 2}|l  ��P������h�	hd"����DEFSCH [R|�Q�<��b�@Default Schg���n� ���������� K"4�Xj��������
)�FB�KLOG1 @z��T�῀  U gy��12=O�����5LG_?CNT  �����)�IOEX 2ڱ����A ��C��]$@������!��
Weld S�pee%��IPM  d$�/�/�/�/�??(?:?��OTF 2��A?�?��?�?�?�?C8=�����@����?K)�PCR 2��p&I�BH�?��BC!�FK<D7������?�ffAZ �A"��OjFM"@���㨶/�O@O"@������WOELG���k%*_�F�023�45678901JRUK%4_y_�_�_HI�ȩ_7]�OOSRA%M2��IB�$�_o�CRGSEL R�<�Q� 	P�rocess 1HoSf2�_oj3iU�o4i�o5�-(mlXS���o7��kn�8i'l"@���� �_);Es-B� �W�%V�oltage�2�qsfc%Dw|!�@]y�h��a�Wire f6�  s�$	� h c%[&t/�oDS�l*� <�N�`�r��������� ̏ޏ����&�]+zv�d"����  �#��E�Z"!��a���^/�� ��V𾔩a�aɒCu�rrent�Amp�=���l�eu� ��Q�c�u��������� ϯ����)�;�M� �W���a�����ឱ	q ��)q��Iq��R�͹� �g�a�aA��b-���-�@	q-�)q-�VE!��\�e�	q?�����Z�%������ϻ�������PDRuS R\zH��jq��C�U�g�����gߩ߻�u� �ߙ���������]� o�)�;�M������ ���#������k�}� 7�I�[����������� 1C��I�� Wi������ ?Q/��� ���//)/;/M+ �U/g){/�/�/M/�/(?cS2�S^=R���b�S2UPYp^=��=�o?�33�H1>E0=L��>TI0h!�"�#�1$�1t9�g�q�#�?�v�#>�8�8CW�IRE 2&M<��?�?h�>�3��>�G(=�J*��ESCFG ��G�A��Y��OOˎE�7])COUPL�0
=k
0�vkB`�D �^�L�[�OZW�O�G_��OP_G_Y\�HNB � ��Ec&FUST_OM  =k
8���y�O&EEMGOF�F !=kS��~)BPCR "�_&�@���zqC{sU� �MJo�\zt�f_oeo��
Cl�q¨1