��   	��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����AW_SCH_�T   � �$CMD_VOL�TS  6W�F?AMP?PK�U
FREQYUL�SE@SPEED�@TIM�FDB�K:�UOMME�NT ���$$CLASS ? ���������� VERS�ION��  ���IR�TUAL��AW�E*  R �� t $ <�A�  +��?���F�����FX j|������ �//0/B/T/f/x/ �/�/�/�/�/�/�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�O�O �O�O�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� �������� *�<�N�`�r�������Runin�����م=��ͩ�	� Burnbac�k��
��  W?iresti2���@����ٍe� On?TheFly?�