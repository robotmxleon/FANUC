��   ?Q�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����MN_MCR_�TABLE  � � $MAC�RO_NAME �%$PROG�@EPT_IND�EX  $O�PEN_IDaA�SSIGN_TY�PD  qk$�MON_NO}PREV_SUBy �a $USER_�WORK���_L� MS�*RTN�  �&SO�P_T  �� $�EMGO���RESET��MOT|�HOQLl��12��STAR PDIU8G9GAGBG�C�TPDS�R�EL�&U� 9�� �EST����SFSP�C����C�C�N	B��S)*$8*$U3%)4%)5%)6%)�7%)S�PNST�Rz�"D�  �$�$CLr   �����!������ VERSION��(  ����!IRTUA�L�/�!;LDUI_MT  ��� ����4MAXDSRI� ��5
4�.1 �%� � d% ��}? i?�?���" ���?�?�? O�?�? 6O�?3OlOO-O�OQO �OuO�O�O_�O2_�O �Oh__�_;_M_�_�_ �_�_�_�_.o�_Roo oMo�oIo�omoo�o �o*�o`� 3E�i���� &��J�������}� ��e�w�쏛����я �X�C�|�+�=���a� ֟����џ�͟B�� �x�'�����]���� �����ɯ>��;�t� #�5���Y�ο}���� ��:����p�ϔ� C�UϏ����� ߯��� 6���Z�	��Uߢ�Q� ��u߇��߫� �2��� �h���;�M���q� ������.���R�� ���������m���� ������`K� 3E�i���� &�J��/� �e���/�� F/�C/|/+/=/�/a/ �/�/�/??	?B?�/ ?x?'?�?K?]?�?�? �?O�?�?>O�?bOO #O]O�OYO�O}O�O_ �O(_:_�O#_p__�_ C_U_�_y_�_ o�_�_ 6o�_Zo	oo�o�o�o �ouo�o�o�o �o�o hS�;M�q ����.��R�� ���7�����m���� ���ǏُN���K��� 3�E���i�ޟ����� &��J������/��� S�e����ׯ���ѯ F���j��+�e���a� ֿ����ϻ�0�B�� +�x�'Ϝ�K�]��ρ� ��߷���>���b�� #ߘߪߕ���}ߏ�� ��(�����#�p�[�� C�U���y������� 6���Z�	����?��� ��u������� ���� VS�;M�q ���.R �7�[m�� �/��N/�r/!/ 3/m/�/i/�/�/�/? �/8?J?�/3?�?/?�? S?e?�?�?�?O�?�? FO�?jOO+O�O�O�O �O�O�O_�O0_�O�O +_x_c_�_K_]_�_�_ �_�_�_�_>o�_boo #o�oGo�o�o}o�o �o(�o�o^[� CU�y���$� 6�!�Z�	����?��� c�u������ �Ϗ� V��z�)�;�u�q� 柕����˟@�R�� ;���7���[�m�⯑� ߯�ǯٯN���r�!� 3�������޿����� ÿ8����3π�kϤ� S�e��ω��ϭϿ����F���j��+�
Se�nd Event�s�S�SENDEgVNT��Q����� %	��Datya�߶�DATA���ځ��%��Sy�sVar;��SY�SVw��ڗO�%�Get�x�GE�T+��%R�equest M�enu���REQOMENU?��ۚ� ]ߞ�Y���}�+����� .��d�7 I�m����* �N����� i{��/��/ \/G/�///A/�/e/�/ �/�/�/"?�/F?�/? |?+?�?�?a?�?�?�? O�?�?BO�??OxO'O 9O�O]O�O�O�O__ _>_�O�Ot_#_�_G_ Y_�_�_�_o�_�_:o �_^oooYo�oUo�o yo�o �o$6�o l�?Q�u� ���2��V��� ������q������� �ˏݏ�d�O���7� I���m�⟑���ݟ*� ٟN������3����� i���𯟯�ïկJ� ��G���/�A���e�ڿ �����"��F���� |�+Ϡ�O�aϛ����� ߻���B���f��'��a߮�]��߁ߓ��$�MACRO_MA�XX�������Ж�SOP�ENBL ���2��ݐѐ��_���"�PDIMS�K�2�<�w�S�U���TPDSB�EX  K��U)�2�����-�