��   K�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_���$$C�LASS  ������D��D�VERSION�  ���/IRTUA�L-9LOOR� G��DD<x$p?�������k,  1 <DwX< y�����C�����	/��Z�Zm//��/_/�/�/�/$ ��/�/	?';�$M�NU>A\"� 
 <��4/d?��[=�-/�;�i� CI��?�?�;DD@#�c���?�?{9@ 'v@ CF�3O�?[O�= cO�OwO �O�O�O�O�O_�O_�E_�;5NUM  u���� tU�TOOLC?\ �
Y?O�_Cj�� GO�_	o�?o?o%o7o Yo�omo�o�o1_�o�o �o�o;!CqW y�����sV�Q �Vy�Wy