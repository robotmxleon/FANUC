��  U��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A0  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ����AIO_CN�V� l� RA�C�LO�MOD�_TYP@FIR��HAL�>#INw_OU�FAC� �gINTERCEmPfBI�IZ@�!LRM_REC�O"  � AL]M�"ENB���&sON�!� MDG/� 0 $DEBUG1A�"d�$�3AO� ."��!_�IF� P �$ENABL@�C#� P dC#U5K��!MA�B �"�
f� OG�f d PCOUPLE, �  $�!PP=_D0CES0�!e8�1�!  R1> Q�� � $S�OFT�T_ID�q2TOTAL_E�Q� $�0�0NO��2U SPI_IN�DE]�5Xq2SC�REEN_NAM�� e2SIGN��0e?w;�0PK_�FI0	$T�HKY#GPANE��4 � DUMM�Y1dJD�!UE4�RA!RG1R� � $TIT1d ��� �Dd�D� ��Di@�D5�F6�F7*�F8�F9�G0�G�G@PA�E�GhA�E�G1�G( �F�G1�G2�B!�SBN_CF�!'	 8� !J� ; �
2L A_CMNT��$FLAGS]�CHE"� � �ELLSETUP� 
� $HO�ME_ PR<0}%�SMACRO�ROREPR�XD0D+��0��R{�T UT�OB U��0 9DEVIMC�CTI�0�� ��013�`B�Se#V�AL�#ISP_UsNI�U`_DODf<7{iFR_F�0K%�D13��1c�C_�WAqda�jOFFu_U0N�DEL�h�LF0EaA�a7b?1?a�`$C?��PAb#E�C#sATB�d�� W_PL�0C�H/ <� PUD�P�B
2ds�`Qg�dsDUT�PHA�gpSF���WE�LDH2/0 �=Lc7w7atAING�0$�r�1�@D2�4�%$AS_LIN�;tE�w�t_��2U�CC_AS
BFA�IL�DSB"�F3AL0�AB�0�NRDY��P�z�$�YN�Wq<��`DE6r��`���+�����tSTK��+�;s7�;sNO�p��[�̈́r��U* Ȁ%�9 �  �� ��q`�G�C�G�+�U�S_FT�vpF��ǂG�SSF��PA3US���ON7xǓ�HOU�ŕMI8�0�0ƔSEC�2�r2yi �rHEK0�v�8vGAP�+�	�I�� � GTH���D_I���T= �l� ����`�s9!̅����9!G�UN1���q����#MO� �cE 	� [M�c�����REV�B7�� � �AXI� �R�  � OD��P-��dPM��!%�;�/ �"8�� F�q�P��0}DfT p E �RD_E%�Iq$�FSSB�&$CHkKB�pEdeAG� ��p�  "
�Ա� V�t:5���3!�a_�EDu � � C2��qS�`�vl ��d$OP�0�2��a<�_OK��Y�TP_C� <�d�vU �PLAC�^}��p<� xaCOMM� �rD|ƒ��0�`�KO]B�� BIGALLO�W� (K�w�0VAR��d!�1B �P0BL�0S � !,K|aԚPS�`�0�M_O]=՗��CCG�`N�!3 �� ��_I_���� �0�� B.��1S|� ~�CCBDD�!��I�����@��84_ �CCWp�` OOL�
��P'�MM
�n�CHs$MEAdP�d`qT�P�!��TRQ�a��CN���FSa3��ir�!/0_F��`( D�!�� CFfT7 X0GRV0�z�MCqNFLI���0UJ�����!� GSWIl�&"D�N�P��d��pM� w� �0EED��@!��wPo��`�PJedV
�&$�p�1``�P|��ELBOF�  �=��=�p/0���3!P�� ��V�F����G� �A0WARNM�`ju��wP��8�𼠤 COR-��8`FLTRjuTR�AT Tlp� $7ACC�rTB� ��>r$ORI�.&���RT�P�pg
`C�HG@I��3�TH{�1�I �r19K��� ����"�Q���HD���a��2
BJ{PC��3��4�5�6�7j�8�9�COfS_rt���3��V�OLLEC�>�"MULTI�b
2`��A
1��0T_�R�  4� STQY2�R���).���p��o� |�A06Kb�Ib$��0�Pc���UTO=�cE�EXT!Y��
B!�Q 2 )
l��a0��R�u�r����   �"���Q����qc�~#!|��1Y�qM
�P8$  l�TR�� " L@q��/��P��`AX$JOB׍���:�pGx# d��? %?78��3�p%��~�CO_MOR��$ t��FN�
CN9G&AF�TBA�� �6�JC��9��D@r�.�1CUR.KPa`/E,�2��%��?��t�taoA��XbJ��_R��|rC�LJ�r�H�LJ�DA���I������2G�� �C}RfT&� ���bG���HA;NC6$LG��iq da��N�*�YaCᇁ�0T|rf�R'L��mT�X���nSDBWnSRA�SnSAZ`�X��8$  ' FCT��e�K_F��Pn�e�M
P
�QIkOh����� �1��e���Cg���A���MPa� ��HK�&AEUp�p�Q����9 �'  �]PI��CSX9C��Zq( xs��sR��T�R�CcPN��v��MG�IGH"���aWIDR�$V�T�P��9�EF�P4A cI�XP,aQ�1u�CUST��U:��)R"TIT���ڋ%nAIO�����P_�L���* 1\0��OR��$! �q���-��OeP�� jЅpIp�Q�u�J8��
��0��DBPX�WORK��+��$SK0���T�DB�T)PTRw� , �l@Ab��s�R0�bؠD��A:0_C��0��=�+`H�PL�q��"R�A�"��#�D��r�B����BJ���9��6� jDB�Q��-�r~qPR��ΰ
�
�Dct��. ��E�S�a���L2Ӊ/��b�@�( ���0�R�Pj� Y1%�b��A�E���� 2D�7���R�E���3HPC~�  .$L���/$Ӄ�����IN�E׶�q_D����ROS��E0"2q��f0�p��PAZ�tAsb�ETURN����MeRQ2UR@�CRŐ�EWMwp��SIG%N�A&rlPA��W��`0$Pfg1$P�P� 2j�B��q����!��DQ���f������׶GO_AW;0���vp���qax CS'���C%Yx42O�1�8�T8���2��2�N��@��CtDۣDEVI�ѐ 5 P M$RBֳ��I�yP.�i�I_BY��q���T�A9�HNDG�6�������b�DSBLr3ͳ��7�Le7 H� �� ��TOFB̶�FEБg')�h�ۣ�f8��DO�a�� MC9�"�`�s(r�(��H�PWp�N7�SLA4���9IINP!Ѐ� ж�ۡ��:D *�S PNp�#�lƍ�1��W�I1��J��E�q�87�qW��NTV�#��V ��SKI�STE^��b��pڥ&�aJ_�Sjb_>����SAF�k���_S}VBEXCLU�*�po�D�pLX ���YH��%q��I_V<9`�bPPLYj���p�����_ML��}L�VRFY_D��M�IO�`  P�%`�b�Oe��LQS�|b��4}������P�u���6Y�AU NFzf�� ���)��#�cD�4Ͱ�� S��r�AF� C�PX����&`� ;j��pTA#��� � ςi�SGN��<��<@3�P��c_� t�a���qd��rt��`UN>�����<@rD�p]�T`����%`������p�pI>�= �@��F��\tG@OT S����|������塁�@y Mr�NIC>�2K�GM A��iD{AY�sLOAD�虄D��5�� �E�F pXI�?j�ď�~cO� �5�_RwTRQU�@ D��t��0Q�p �!EԠ��< ?K�%�>`� �M�AMP*Pp��A�"'; DB�'��VDUS�U�.�CABU�B`��NS9@ID�1W�R$�Q!`V[�Vq_#< ; �DI@�J$C� /$VS�SE�#T�BDC�A�� ���|�DB�AE_l�;VE�P�0SW!�!�@x�3�2� @�`�OH�@3PP <IRwqDBB�p�=�!U����t"BAS��o'~P�Pn%[�d� B	� ����RQDW]%MS�� �%AXC'�;LIFEC���� ��	2�N1EB5��3EBChd@/Ź�Cq`ʡaN�4q�6��OVՐ�%6HEh�DBSUP$�1��	2D�_�4j�BH1_!C�5š�7Z�:W�:qa�7�S��"BcXZ�PʁEAY2HEC��T�pސ�NM��� �q0P�dD �`L��@HE�VXCSCIZ?6k0��[�Nh�oUFFI�0�� C��������6��zrwMSWJEE 8��KEYIMAG�TM���S�A5��F��|
q�BOCVIE N�qF 	�PLQ�_��?�@@|p&`KD�G� ��ST��!>R|�FT��FTD FT|� FPEMAILb ��aA���FAU�LSHR�*�;pC#OU_��q|pT��U�?I< $�S_��S#�ITճBU�FkG�kG@�jp`p�0B�Tk�C��Rws�PSAV(e�R�@+Bd�$ Cg�p��P/d_ň�$̰_�Pec F�iOT����P@�0���jA�gAX�sq�:p�P��\c_G3
N�pYN_e!�pJ0QDf�W�r�d"MO�_0T��F��
C�E2���^ЈqK��ey&^�5q�)�4��qL���nq�S�cC_ܐ��K씐pu�t��R�A�u�XnqD�SP�FnrPC�{I�M5c�s�q�nq�U`�w{0�0��PIPR�dnsN!DB@�sTH���"ûr� Tߑ�sHS{DI�vABSC_�9@`�V��x�v��c~�,���NV��G��~�H*@�v�PF!�`d�s0p�a��SC�\��s�MER��nqFBC3MP��mpET�⌐mM�BFU�0DU�P0?�M�B
�CD�yH�l�`�S��NO��
��N� %�i�cg�V�PSf�CB@v�	C���aBAd��`U OH����c d�� �����}�锍��9��D疢疮A�7
�8�9�0��U1��1
�1�1$�U11�1>�1K�1X��2f�2���2
�2��2$�21�2>�2�K�2X�3f�3�3T��
�3�3$�31�U3>�3K�3X�4f��jrXT�TP < sK�p<6p�p2Ǻ��C@FDR�QT�PV��b	2�p�v�	2REM�F���0BOVM�s��Aޟ�TROV��DTl3`��MX��IN��8Q0�ʶIND����
	�i��`$DG@�a{#��4P5�D����RIV"�=20BG�EAR�qIO�K��;N0p}ة�(����@�0<Z_MCM�@	1�F|0UR�"�R ,t� a?3 P0�?��!?��EG��*QHa��e�S� � P�a��RIM�P�SE�TUP2_ T D �STD6���<������I�C�Q�RBACrU T[ �RTt�)Nz%��+p�IFIQ!+p��А���PT{b�&�LU�I1TV � Y�PUR�!�W2�r�<qv��P�� I��$��S��?x#�J�QpCOw`�cVRT|� x$SHO���SASSY��a?5�8�
���A�W��RFU��15q��2pfu��*@�X |�wNAV�`���3���*@�R=1��VI3SIJД�SC��遡E�c�\�AV��O*��B%EX�$PO��I\ �FMR2b�Y o�X�} p�bpNt�{ߍߟ߶�(�P���_f�G�_��B��M4�Y�k��DGCLFR%DG�DYLD��7�5�!6.�04\�MR�3SZ��P�	 T�F9S�`2T[ P!��|bs�`$EX_����1�`Ā\2�3��5��G��9\R��
���PWeO�&DEBUG��"���GRR�spU�BK�U�O1�� 0PO� ;)' ��:' Mb�LOO�ci!�SM� E7bA ����� _E ]� �@h� �TE�RM�%^�%��OR�IBq� _�&C@SM_OpL� `�)���(�a�%*QUPRbg� -���]�#0^��G:0E�LTO{Q$US]E��NFIc1G2���!���$4_$U;FR��$j�A1�}0=�� OT�7��TqAX�p��3NSTCp�PATM�d@�2PTHJ�;�E4P_bD�H2ARTP`R5�PPa�{RG1REL�:�aS�HFT?�H1�1�8_�N�R�8��& � $�'H@a�q�B���b�SHI@�U�� JaAYLO��a�a����Y�1��~�J�ERVA�3H7�Cp�2�����E����RyC�~�ASYM.q�~�H1WJ[7��E ��1Y�>�U2TCp �a�5�Q=��5P��@,��bFORCpMK%�GRz!:c��'"`&��0w0�aG_�HOb�fd Ԟ2��& �X�OCA1E!��$OP����V�t F����P��P��2`RŃ�aOUx��3e��R�5Ie h�1���e$PWRL�IM;e�BR_�S�4��� �3H1UD����Q�Bte7�$HSu!^�`ADDR2�H}!G�2�a�a�alp_p��.x�f H!�S��񀌳u��u
�u�SaEv��h�2 HSH��:g $���P_�D�H Y�RrPRM�_��^HTTPu_i�Hx�h (*��OBJ���b��$�2�LE�3�s�i� � #�"�AB%_
�Tp#�rS�Px����KRL{iHITWCOUw�B6�L `�rQ��U�`��`�SS��JQUE?RY_FLAQ1�pQWR�N1x�jpgP&��PU����O���q��!t��/t��� _�IOLNw�k(��� CJq$SL�L$INPUTM_Y$;`��P,���̀SLA� l׀�(�$��C����B��IOgpF_�AShm}�$L ��w��8AِU� 4@�_1��݃��情@HYp1ǧ���W�UOPen `l�ő2��������[`P�c;`嗠	������2Ja�oo � K�NEaG�4�v7F�Da��2J7zVpOQR$J8q��7�I_1z���7_LAB�1�P|���p�oAPHI��Q{�:��D�J7J�-�ީ_KEY� ��K��LMONzx�p�$XR_����)�WATCH_p��C��D�ELD��1y�P��eq @Р1qV�@&�U�CTRC�U�i����LG��ro� !#�LG�Z�Rࢵc��c���FD��I����\!�� ��� ����e�Dqf�c e�c�e�ΰe�� e���@0J_�ѐ1j��qʦ�F�AxǒĞ�Cd9(��SB����@c��c���ΰ��I������ƍ �ƞ�RS���0  (_L)Ne�<sѐ�� �)��6Ѽ�UosD�r�PLM�C�DAUiՃEAwp���T�u�GqH�RNqo�BOOw�t� C���`I�T\���� ������ScCR���㇑DI��Sw0HRGX �� �z�d(��o���w��W�o�X�z�JGM�^�MNCHl�n�F�N�a�K��PRGƅ�UF��B��FW�D��HL��STP���V�� ��Г�RES�HzP��w�CdD@��1Rz�: :�^�Unq���9���H�k�����G w�@( w�������s�f}�OC/ ��EXv��TUI��I��7� C�O�����<@����	$��<@��NOANAo�A2� gVAI���tCL~UDCS_HI$��!s�O�
�S�I��S��IGAN���ɳ��h�Tcn�DEV<�LL�ALʀo�BUI �uP��j@T��$��E�Mr���]�.+!	1vP�j@ހ��~p����1�2�3����� 
0w �C��x�Qp@5������IDXa$�9 [����֥1�ST�ƐR��Y� <@   _v$E.&C.+��pmp=&P&�!��	1x L����`��4@r�`Na�eENwp�d0�?���_ y �ap7�}p	b���#�{MC7�z �C��CLDPƐUTRQLI��TT�94FLG)"0�Q53�1DD�57t�LD55455ORGT�8�H2_� �F�8!s�D/r �#�S?{ � 	59��455S�PT0���0y0�4�6RCLMCD�?�?Iƀ�1��PM�p^���|�?$DEBUGGugQODATAY��T ��UFE��T)!���MI6p�T} d�@��RQ��0DgSTB�`� �F��HAXR��G�LEXCES$Rh!�B)MZ`��~���B4PNq�BSq�����F_z@�H�S[�O�H�0wJPTH�� &P�v�m��QMIR� �� � []�R�RCT��N}���VO�ZA�ZL�RC��PC��Q�`D��O��^�CURPX+_THqG�P�`R` |1h )`/d55R^`�`yS�P �B_FR@^�a\fZ_��^ddp�G��* TP�MK�H�� \��r�Fv$�MBu�LI�q�cR�EQUIREG�M�O�lO�kfB-��1L:� MG�� ap����`|��cB�MNDU�Sz�>�5�Z�29sD��Q�IN�p��Q�RSMf�Sx� �Q��!E]�qQ'qP�ST� � 4f�LO�P�RI �v�EX�vANG�X�A��1�AQG���@c$�QG��MFh� �����"��%&�2�N�fSUP�%�!F `�RIGG�� � ��0�#1��Ӫ#Q��$$���%#n�א~��א��rP��wAZw@ECTI9�~��!2�M\pn9� t�pMD�I��)��� �DA�qH�pu��DIA���ANSW,��wT���D��)RAO7�\�0�Љ �QU���VB�70�A�AO�_V@�ъ �C���sLX@�b|ٰ��P��h�v���P��KES�!���-$B����� �ND2FB��2_{TX�$XTRA�41����`LO�Ъ�1�$RG��B F�8��|�g�_��QRR2>�E�0 #W�e��A�1 d$CA�LI�@2�G���2��RIN����<$R��SW0"DᣫwABC�xD_J���a����_J3�
��1SPs�rp��P��-�3,���?���B\�J�l��2�1O8�IM� �2CSKP ":��~�YÛ�J���2�Q��̵��̵·�p_cAZ�2h���EL<g�FAOCMP�s�1�!I�RT�A)�Y�11�i�G��1�K�> :Y�ZW�SMG�܀v�4JG� SCLP�uSPH_� �0���������RTE�Rࠧ�P�IN��ACz�|��� ⲼA ��} _N�я�������1���?R�� �DI��0i DH�P3��ё�$V0��Rs��>$v��pP�1����@Ro���ВH �$B�EL�?w��_ACCEL��ث�Ц�P_Rـ� �QT�!�*aEX2L 6b��3���׀c��.aУ����36cRO
Q_�m�J�P��2�p�`��_MG�$�DDm�����$FW�0݀�Ӊ�Ӥ�~��DE��PPABN6��RO��EE`� ��0±�YAOP��h �a_��YPaPCD��YY����1 �!YN�@A��7�����7�M�A��ig�OL�de�INCa��q������B�����AENCS��Á�B�Ѥ��D+`IN"I6b��ހ�ďNTVEk���2�3_U�����LOWL�#F�0��DF�D�`��� ��r`RC����MOS� �wT�PP�2��3PER/CH  8OO`�� z�q�!�4! $��!�)b��A6b�L�tW����F�
�4TRK��!AY[�(cOQI6bXM��p/�SQ�� MOM c��BOR�0���D�㣧ad��⍠DU���7bS_BCKLSH_C6b��@YO`�?����*N�ĵCLALM���1�?P�6%CHK0� �GLRTY������Ѕ�|1܁_�N_UMzC�&CzC{���#��7LMT)�_L�0��$+��'E�-� �+�  ���%��>��C�!4�PC��HI��`q�%C@8�{��CN�_��N"C�6��SF�ѯ	V!�p!����U1���5Y8CAT�.SH�����?a���`X�7aX�L�n�PA�$&��_P�%s_����@Pn ��`rDc%JAa�PfC	 OGs7�TORQU�A�Li����bd����B_W �IU�n��D_��EeӪ�EI�KI[Ie�F��P�As�JX��w�VC"��0�jS1q^o�8�_��wVJRKq\�R,�VDB��M���MPp_DL_��GRV�D�T_��Te��Q�H_^��S�#jCO1S0k1�0hLN�PSk tUZd_�Uiv�Ui'Q�j�lEQ�UZN`d�QM�Y\a�h<b��Dk�iT�HET0$NK2a3e�rY�]`CBvkCBY�C��ASrq�Dr'TRq_�RqvSB8_�pr*uGTSֱ��C0��qO�;C_Ǧz�c$DU` ��r�� ��xR�v���Q��53&�NE��7�I^`q#$;��$=�qAu;�pD�"e-h-aLPH0e����StU��e����e��f�����f=�V�]�VR�O�u�V��V���V��V��V��V
ɋV׉H]���|�t���1����H��H��H���HɋH׉ON�OR]�O�s�O��O��UO��O��O��OɋO�fF�?q��e���P�SPBALAN�CEc�=1LE�pH_uSP��pf�f|�fPFULC��`����e��1�+��UTO_[ �ET13T2_���2NB!�� ������ ��p�Қӊ�T
O����@I�NSEG��=REqV��= ��DIF3f�1��1�1�&COB�&!�S�2�@���M!�TLCHWA�R��&�ABBA�$MECHHq�`V�,\�q&AXVP4u�84�@�T�� 
v��A�b���ROBn CR����j2 �M�SK_֠�ԓ P+ j�_�R���2����51�2���������$��>�INű��MTCOM_C|\P�Д  h����$NORE���Q��.�@�� �4�@GR�Ba�FL�Aű$XYZ_�DAQ����DEB�U��Pf�.�mЖ ��$/�COD!� �҇b���$BUFINDX�������MOR��� H�����E&���~�^�$޲��Xo1�� TA��� ��ѰG�Ҙ � $SIMULp@�С��\��OBJ�E��\�ADJUS<z�m�AY_I�A�D��OUT�@�Ԡn_�_FIb�=��T�@��������q���������D,�F�RI��T�RO�@��E�A�OPsWO�P���,�ПSYSBU+���$�SOPT���;!_�U<^��PRUN0҅�PA��D��`�Y� a_��2z��AB���
0��IMAG!4���PϱIM����IN�P����RGO�VRD�v�e��P0����� ��L_R�zA�(�"�0RB� � >1MC_ED��b� 
0N+�MW	1��MY191��SL����� �ޡ�OVSL��SDI5�DEX�3��3$
�V�@�N��A���� ���n�C��0T����_�SET�@��� @0�@!��RI^����7_Lq@YL���x�0 ���Ta��@ATU}S�$TRC�8��ҔBTM��	I��l41sU ��� D��E���4�E���� & �EXE�r!L� "��)�0���UPؒ�!IS��XN�N��1ldQ� ��PG>՟L�$S�UB��V�ZJ_MPWAI�0P���%LO� ��̰[��$RCVFAIL#_C�i�!R��iЀr�e1�0�4���%�`R�_PLZDBTB8�A�2i�BWD�&Y�3UM�@�$IG�������0TNL�0�$@2�R'�T�~@�@��PP�EED5 �3HADCOW�@c�Y�f�E���4�p!DEFSP>�� � L��|��0_�0���3UNI�����0C!R L��`̰P��@�P1�����Ю@^Ѡ��� ���X�N�K�ETB�@��	@P|42��� h �pSIZE���������`ASx�ORZFO�RMATK�*4COX~ \AǲEMn�|D��3UXC��CBLI�%2��� $I�OM�P_SWI/��E҉�Wi�Js��AX�
0%0AL_ ���@�0"�gPBJDpC��D��$E!��J3D�H� TV@PDCKC m�X�CO_J3r�RQR�Ģ�	_]R��@C�_/1A  � ��h�PAY�qҧT_e1�Z2�S�@J3�p��[�U�V�S6�TIA�4�Y5�Y6�MOM�c$cc$cc;�B� ADcHfcHf6cPUSpNR)due�cueb=��B�ħ?` I$PI��U lq�U*s�Uus�Ujs�U Ut�f�kit�t��v��v_!��m���:v3HIG�Cv3�%�4iv �4�%� ��iv�sxx�!8�y�!�%SAM���p�tiw�s�%MOV��$�'�
�ް)p%�� � #��0�P2��P%�0� 5�`!��@��H��#�INj��@�sq���h���"s�������ӋGA�MMǦ���$G#ET���Є�D�T/�=
z�LIBR9!W2]I��$HI8 _��H�%�H�E"�U�AO�r�c�LWJ�����r�@��c��Rn�M0�AC5x0� a ?^I_�p2�/��B�X�A�Y��$c/�Hf��C ��$,X 1U���IXRk�D�0>�A!�$@�LE �8q�`���Xq��Z0MS�WFL�$M�@SCRI(7���)q�T"p�0�A����P���UR�$�v�KS_?SAVE_D-B�;#NO�PC`<"�T B�&��_�a�YW��i�Y �`����pkR#uܸ�SD��p#�s0�@�,� $�cxY�svY�x@�<Š���<!p�@M�ũo � "�YL�c��Y��S��6�0 �� 0����J�������H�	�t�Wq�����`��1�t�M����CAL���Q��o �1T"�@M3�*� � s$��G$WR� �����QR�oTP�vT P�}TP�T0���+�(�C;�@X�0O~S�A�Z�տ@��Uԫ �ՑOMK��V����p����̿`CON��N ���@�Q_v"� |=Q�B�$i�� c��cB��Z���j��A �D���t�P��P_A�PM� �QU�p � 8�@QCOUM�i�Q�TH/0HO��G�H�YS�@ES�F�U�E2�8�E@O�D� � �@P0�@�`UN�����0OVr�а P����%$��W2�ROGRA���22�O����IT�����t�INFOXѱ ��A����ȩ1O�I� ((�SLEQZv/Nu/ �����OS��s$� 4�@ENAB~�� PTIONZ�4(r�\�4cGCFl�0�J� �A���,�R�����OS_sED� �е �NR��K�:G�E��sNUAUT^�COPY�8 7�1j�MN�NAEPRUTf� HNֲ OU�Bo RG�ADJXѶTBX_t��2$�0��мW�P����v3���#EX� YC~�^{�RGNSh����ޠLGO��PNY�Q_FREQ�bW`��MvM!�D��LA���D!�c��@CRE�3�R���IF�a��NmA�q%�$_G}4�TATB0�$>�MAIL�r2��!��B��1x�!1�$ELEMl� �s0vFEASIy@��L���2@@K�66�V�2�I���0�D"8qJ��k2AIB�APE��vpV�!�6BAS&R�52��aqU�p��W�$�1~�7RMS_TRe3 �A���3�ӓp�r�!�4c N�!"������	B2 2�  ���ԇ�(F�2'G�2/��_����2SG�g��DO�U��N�!"PR�e�m �6GRID���b�BARSZwTuYz �OTO?`�Xѻ ��_�$!���B�DO��i� � ����PORp���C�f�BSRV� Y)TVDI`�T�P@0QCT� MWCpMW4KYU5KY6KY7KY8/Q�)�F�l��$VALU�35�(42��r�Fh�� uY����C�!2�� #AN4��R�!RR!>2�TOTAL�s�a�2cPW:#I�AHdR�EGENFj[b��X��8��R%��V-�TR�3�rFa_S8��g[`��V���b��2E��#�@L�1�-cV_H�@DA-��`pGS_Yf���^&S�{AR-�2� �IG_SEC�`R2�%_���dC_�F�Q��E�q�OG6�kjxSSLGEpl�� >� _%��/�0`9`S���$�DE.QU>����sT�E���P�� !��a��aJ�v^�3IL_Mm$;����`��TQ-�6���0Ƨ��Vh�Cv�P�#1��mM��V1��V1��U2��2��3��3��4��4��$��`ӓ%��� 0����INA�V�IB=�p�]��d�2�`�2l�3`�3l�4B`�4l�X�WB�SB�����D $MgC_FP���%��LC�B�f#cMo�I��oC ��6��q�L�KEEP_H/NADD�!#��0-�C�ѫ C��A���D�O&�"�{��3�pD��!a#D�REM[��C�8a�B������U��$eC�HPWD � #�SBMS�K�BCOLLAB�/��P@�$a�" I�T$ ��fȕ��� �,(�FL{�W�M�Y�Nڐ1�M��C`r�~G`UP_DLYX�=��DELAc�9aZ�"Y�AD-��A�QSKIPw�� i�P��O��NT9�����P_����� �ҏ�÷�aѹ�ѹdP кqPк~Pк�Pк�P�к�Pк9��J2�R ���qX�0T G#r���qr�� �r�����)�RDCS��+ �_�R�R1�o��I�R�!��J��*DR�GE� T3�ÆBFL�G'����*DSPC���!UM_r�!�2/TH2NrA<�e�� 1� ��E�F� 11��� l`����O�v�ATy� �.��Q&������� � *D�Ҙ�I�H���W U�2]��c�`u߇ߙ߽߫� T�3]��������(�:�L�4]��]�o��P����L�5]����@�����"�4�L�6]��W�i�{��������
V�7]��������
\. �U�8]��Qcu������S�L�  ��1V�p`ДUЙ�E%$рp�e)f&cIO��Ip�W�R��WEC��# M0����#d� �+��$DSAB] � �""c^�CB�,p_�RM
E�+��	�D��0E�"��M�D"'�!�D� D��p�'DBG_~@P0D�3%!eaPG
A@���ա�S232Ni� ����P��pICEU�2!`k$��pARITq!aO�PB�rFLOW>pTR(.b��@q�CU� M%3UXT�A�qINTER�FAC�$��U`���SCHA� �t�ݐ"!hp�$L�`�`OM'p�sA��"�0Iᓴ0Q@A+Ӫ	TDSv`���8c3�EFA����r��S� k��`8b �q��R H��6A �ٶ�q  2� ��S��M �	�' �$)�s�0�
e�C2`_%pFDSP�)FJOG�`�#�p_P���"ONg�u����'�	6Ky0_MIR�EAb$wpMTY��CA�PK�wp4Ц@�4"AS�p}@r"At �EBR�KH<16=��R�� �B�s�BBPo0�bC�@BSOCF��N�UD1pY16���$SVi�DE_O�PGtFSPD_OKVR�k��DTR&WCORbW� N�PcV�F�@�WB@OVEES!F�Z^p�S,rF�V t�'�UFRA�ZTO��$LCHa�u�2�OVST��B@WQ���BC�Z� r&PQ@]s  �@�TIN�``!/$OFSC`C�0@�WD|QdxQ%Q��E�?PTR�!e"�AFyD���AMB_C�
�bB5@B<��!q�b�a�cSV��L�k0��ds��RG�g�HAMt�B_=0�e-b_M��`2�:`T$C�A8@�D�B?pHcBKo1~6TqIO�qcu�pqPPAWz��qhy�t{uu�:bDVC_W R#�p1� �p���Q�u���x-s�u3�v3`��{�0p@SQqUR#7@~CAB����,Ӟ`���`�h9�O��`UX~6SUBCPU�O@S����� �dp0ݱ���c�d���?$HW_C]��0ݱrpʆ�� �Ð'�$U��D���ATTRI�0��O@�CYCLw�NEC�A)��CFLTR_2_FI�/��v�LP[KCHKՠo_SCT�CF_�cF_�|��FS��b�CHA��d���8�b�"��RSDU��0Q�3��_T�hY����c� EM"��M"�CT��ݰĀ�����2�DIAG5RAOILAC�sx�M��CLO	P7�/V���b3� H�3��sPR�pMS+� 90��C�qz� 	,cFUNC���1RIN���$0D����!ʰS_"@*?p䣸�Mt���MtGCBLȰ���A�
��
�DA�@�O���LD`0GPpqw�d*A�|�w�TI�����AĀ$CE_gRIA��AF��aPn#ò%`ȵT2d�1C}3�r�aOI�fDF_LY�Rl1�0�LM`#FA  HRgDYO�AM`RG|��Hސ�Q� W��MULSE��3��8P�$J_ZJzR�W�[�FAN_ALML�V�#��WRN��H�ARD�@o6��2$SHADOW ` �����V���!�Q�EY_`s�AU��R��~2TO_SBR���6@(�逺sá@�M/PINF8`��SԜm�^�REG���D�Gy�K�Vm0��FDoAL_N�dFLۅ9�$Mm�l�>g �O`L�K$3$Y("V1�2#��� ��CE!G[CGP
�A ~�/U28S�;��EAX�E,GROB)JREMD)FWR  �A_i�SSY�@D��@��S���WRI  �ɀSAT�*C0�@nPE�A&�w� �"@B���9a��5k�pOTOrn�%`ARY)C`�e���[@FI�@~pC$LINK��GTH2��0T_���9a%�69R[�X�YZo2e�7s�OF�FA`2� \�N�uO	B'@����a� h0��FI���0�?T��AD_J�!�2lR ?�pq������89R� ���	T�AC��FD�UWb$�9x�TURB��X��z!�N�X��� )FL[��PH���� |���309ROa W1�KN@Ms�/U3��{�������W3ORQ�6A����{��@O��N��H�384A��]OVEd("M00J��~��~�Ҁ}F1|J�|�{AN��5�~ȱ)!e}@ ���ve�%�Ә%�6AERSA�	B|�E �`��E$A�Ā��ܥ��V�S�V�AXc�2V��ҁ 4�%8��)b��)w��* �*r�*��*: �*q �*1� �&��)� �)��)��)��)� �)�9�9�'9D1�89DEBU��$�����0��1VbV�AB�V�Tq|Q^VIp�� 
B�s��+E��7G 8Q7Gw�7G�7Gr�7G ��7G:7GqδF Ȳ\4��LAB��)���sGROB�)��2pB_�,&��uS ��%��FQ*U�VAND� |�:$3�_�=!�YW 2qZ�^�mX0�|X5�^�NT��
c�PVEL���QT�~�V�SERVE�PN��� $���A�Q!�PPOHb���`���Q�R�����  $bTREQK�
 ct�
`�g�Ȳ2�e��Q�_ �� l���a��ERR��m"I� �P�NraTOQ��LH�P�$��f�G�U%H��f���b��	a� ,h�Q#e=`��RA�a? 2� d�b{ss�d` ��Ѓ$r����"�eO�CG�p�  >dkCOUNT��`���SFZN_C;FG	a� 4ƀ��;�T�Ŀ���3�����m!��Rs��� �(@M��o���#������uFA���ö�sXd��{�y�a��S��T�O�d�PJ��S�HEL��Yr�� 5k�B_BA�Sf�RSR�֤�"^�S끐�M�1�gM�U2p�3p�4p�5p��6p�7p�8�g@�R�OO��`9�]�NL���LAB�SN�N�A[CKFINpTo����$U��M��� �_cPUV���b�OU�P̠��-��f�����&�TPFWD_KA1Rwa��f`RE�T,�qP/�]��QUE��@�eU �����I���C-�[�[��Py�[�SCEM3A�AAH�A�q7STY�SOސ	�DI�ɠ}s���'���_TM��MANR�QL�[�ENDZ�$KEYSWIT�CH^�s�.�ĔHE�U BEATM��PE�LEvb��@���Ur�F�s�S3�D_O_HOMưO��6�EFA PR��r(v����C��O8�c`�aOV_M�����IOCMG˗?�	�,�HK��� DHX�׍pU�¹�M�x���HFORC���WAR(��R.�OM>� � @�4���U��P3�1��2j��3��4=��Qp*pO��L����b��OUNLO9�����ED��  ��NP�X_ASZr� 0�ЄЍp��$SI=Z��$VAP�e�MULTIP���.�ŰA��� � $H�/����B��S}s�Cr`��FRIFm"pS���������NFO�ODBU ��~P�������U�RN�n��� xU`SI�b�TE�8��SGL*�TA� &opC��C<��+�STMT�\әP��BWe,�S�HOWd�n �SV�7 _G�r� : $�PC�@p7#�!FBZ��P��SPːA�̶� `VD�Оr��� �WaA00 ^T��ɰ��Ӱ��ݰ��T���5��6��7��U8��9��A��B��@���׳A��y���F�ب70���1�1"�1�/�1<�1I�1V�1�c�1p�1}�1��1���1��1��1��2���2�2�2"�2*/�2<�2I�2V�9 T��p�2}�2��2��2��2��2��� `P�>`"�3/�3<�U3I�3V�3c�3p�U3}�3��3��3��U3��3��4k	4�U4�4"�4/�4<�U4I�4V�4c�4p�U4}�4��4��4��U4��4��5k	5�U5�5"�5/�5<�U5I�5V�5c�5p�U5}�5��5��5��U5��5��6k	6�U6�6"�6/�6<�U6I�6V�6c�6p�U6}�6��6��6��U6��6��7k	7�U7�7"�7/�7<�U7I�7V�7c�7p�U7}�7��7��7��e7��7��bVP��=Ub� `{@�e�
wA���Q�U��PR��CM�p�bMb�PR9` ��TQ_+p�R�P�e(a~��SQpY�SL�`�P� � L��jw��A�ؠ; xѠ�D��VALUju�%�x��A6XF�AID�_L��^UHIYZI~��$FILE_L���Ti�$��P�CS�Aq� h ��pVE_BLCK��RE��XD_CPU�YM��YA�us�_�T��B��G�R � � PW-p���6<aLAj�SqAc�RaKdRUN_FLGde@dhaKdv�ke�a@d�aKeHF�Wd�`Kd�+�TBC2�u� � �Bk`(����pĠ���d	�TDCk`|r�b�p��
u�gCTH	�%s�D1vR�~�ESERVE��Rt	�Rt3���`�'p� �X -$}qLEN���t	�}p�)�RA���sLOWI_�Ac1}qvT2�w�MO�Q�S���I�.��B�Q�y�D}p�DyE���LACE,���CCC��B��_M�A2��J� �J�TCVQ�r� �TX�s����������Ѷ� ���J$+���Mۄ~�Jw���R��� ��q2�`������OpJK(�VK��:�>�:�sq/��J0O�>�JJF�JJN�AAL>�t�F��t�n�4o�5/sX�NA1����d�N��DL�p�_Xќ����aC�F6�� `�PGRCOUDPF�Q���N�`�C�� �REQUI9R=rؠEBU��yqn܆$T�2�6��zp ��$$CLA�F� ����5�*�*� O����X�e���~k�IRTUALW��i�AAVM_WR�K 2 ��� 0  G�5a�ͯ٨ʯ.�� ��	��3�*����!�^�E�c���������ɿۿ�㴧�BS�@�� 1�x�� <��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<�~pN�gLMTu�?��7  dQINZl�PPRE_EXEb}� �~AAT��ʖ���IOCNV�Ւ~ �hP�UqS���IO_� w 1��P $����I�4��1��?� ?�`Tfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο�����(�:�Q L�ARMRECOV� �c�L�MDG �(BLM_IF m?����� �+���N�`�r߄ߕ�?, 
 �߾߀9�E�������A�NGTOL  ��
 	 A  � Y�k�Q PPLI�CATION ?��� ����ArcTool� �� 
V9.?00P/03j�+�
88340�����F0����161�2�������7D�C3��+��Non}e+�FRA+�� 6�LP_�ACTIV�	�j��UTOMO�D� �Ո	P_CHGAPONL��� ��OUPLE�D 1� � !3��CUR�EQ 1  UT=	==	�������=_�ARC We=l=�AW�ՕAWTOPK�HKY�Dy�9 'EK]o� �����5/�/ #/A/G/Y/k/}/�/�/ �/�/�/1?�/??=? C?U?g?y?�?�?�?�? �?-O�?	OO9O?OQO cOuO�O�O�O�O�O)_ �O__5_;_M___q_ �_�_�_�_�_%o�_o o1o7oIo[omoo�o �o�o�o!�o�o- 3EWi{��� �����)�/�A� S�e�w���������� ����%�+�=�O�a� s����������ߟ� �!�'�9�K�]�o�����OTOC�����DO_CLEAN��|���NM  H���^�p�������A�_DSPDRYRL���HI��<�@M� �&�8�J�\�nπϒ���϶������ψ�MA�X��������
�X��������PLU�GG����
�PRUC˰B:�H�����d�Oi�Կ��SEGF��� ������:� L��&�8�J�\����LAP������ ���������"�4�F��X�j�|�q�TOTA�L,�U�USENU
���� ߨ���O �RGDISPMM�C� ��C���@@M��O���߹RG_STRI�NG 1��
��M��S���
__ITEM1i  n����� ����'9 K]o�������I/O S�IGNALc�Tryout m�odejInp� Simulat{ednOut-,OVERR = 100mIn cycl!%�nProg A�bor7#n$s�tatus�${ c�ess Faul�t�,Aler�$	�Heartbea��#�Hand Broke���/?�?%?7?I?[?m??��e��w�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O__�?WOR��eKQ �?%_s_�_�_�_�_�_ �_�_oo'o9oKo]o�oo�o�o�o�o�nPOc�!�`c[�o$ 6HZl~��� ����� �2�D�8V�h��bDEV�n�� ����̏ޏ���� &�8�J�\�n����������ȟڟ����PALT�=7�c_�_� q���������˯ݯ� ��%�7�I�[�m��8����%�GRI�e ۱O�����'�9�K� ]�oρϓϥϷ����� �����#�5�G�ɿ��R�=��Yߧ߹��� ������%�7�I�[� m�����������m�PREG;�$�� ��K�]�o��������� ��������#5G�Yk}���$A�RG_KPD ?	�������  	]$�	[�]����� SBN_?CONFIG� ��%!$"CII�_SAVE  ��D;� TCE�LLSETUP �
�
%  OM�E_IO��%MOV_H����REP����UT_OBACKs�	�AFRA:\�� ��^'�`� �<(� �M+@ 2�3/04/01 �14:33:48���/�/�/�/-,��?/?A?S?e?w?�?��?�?�?�? �?�?O�?5OGOYOkO }O�O�O,O�O�O�O�O __�OC_U_g_y_�_��_�_�Ё  (!_�#_\ATBCK�CTL.TMP ?DATE.D:��_�oo,o>o#INI�:�o%7#MESSAGS]a^� >hkODE_D�V�7G�eO���o#P�AUS�a!��� ,,		�� ��ow�o- 9;M�q���������;�����d�`TSK  ��m</Bo UPDT̖`[gd���fXW?ZD_ENB[d3��STAZe�����WEPLSCH �R+   b��.�@�R�d�v� ��������П���� �*�<�N�`�r����������̯ޯ����R�ODނ2��4���/��>� % V�{�������ÿտ翀����/�A�SϾWEROBGRP`���r�GWEWEL �2�D���h��� ��'�9�K�]�o߁���ߥ߷��߼	XIS%UN���D��� 	r����@� +�d�O��s���������METER 92b�_ P��&����J���SCRDC�FG 1�N! �[[?� ������������5/�
QW��M_q�� ��2�%�7I���!GR��Р��o��PNAMoE 	��	$n�_EDY`1s��� 
 �%-�PEDT-v��/*/j�� �����.��µ�����/:����%2�/���/a/ ��G(�//?v/�/?�/�#3g?�/�?�/>�?@�?B?T?�?x?�#43O �?�O�?>\O�OO O�ODO�#5�OoOL_�O >(_�_�O�O�__�#6�_;_o__>�__o �_�_No�_�#7�oo �o+o>�o+ro�o��o�#8c/�//� =��>P�t�#!9/��|���=X��Ï
����@��!CR �/�oG�Y�}"���ԏ��|�
���NO_�DEL��GE_�UNUSE��I�GALLOW 1���   (�*SYSTEM�*��	$SERV�_u�.�G�POSREGP�$r�.�G��NUMu�����P�MU���LAY���.�PMP�ALTǧCYC1�0Ԟ�Ѡծ�ULSUǯ���r����L#�\�BOXO{RIy�CUR_I�~��PMCNVæ�I�10����T�4DLIB@�b�	*PROGRAO�PG_MIծ����ALߵ����B<�G�$FLUI_RESU�(u��j������� ������
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� �������������e��LAL_OU�T 6�q#�W?D_ABOR���i�ITR_RTN�  ����l�N�ONSTO���� ��CCG_CONFIG ��7�7���8�����E?_RIA_I����, ���FCFG �����5_LIM^�2�� �� 	n���<j�ߥ�蜀�dPAV�G�P 1?���-?�C��� C�  CU�b�f�b�f��f�b�f0�DZ`�DD���
�����D�v�DZl~�ʆ��x�D/��9�C�M�Wچa��?���HEp��u�"G_P��1� �� d/v/�/�/�/�/�/�HKPAUSf�16�, ���/ ? 6�?L?2?\?�?h?�? �?�?�?�?�?O�?6O�HO.OlO
O9�?��h�COLLECT_9s	`�N�GEN߰��~��B�A�NDE�Cs����1234567890!W��a�pO_1V��
 H+���)l_�_a�k_}_�_ b��_�_o�_�_	obo -o?oQo�ouo�o�o�o �o�o�o:)� M_q�����h��Fm�K �|N�FIO !
Y �A����������ʏb�[TR� 2"F�(��b}�
�؎��#q�x� %[�_MORm$� �)����� ����ǟ���ٛd��*n%r�, %?	!	!I�>���KH���$�R9&�Ow�v�v�C�4  A��
� �x��AA�Cz � B�fPB���Co  @��������:d�
\�I�S'f�\�T_D[EF*� �%�x+�����INUS��&,@�KEY_TOBL  �,v�� �	
��� !"#$%&�'()*+,-.�/*W:;<=>?�@ABC�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~�������������������������������������������������������������������������������͓���������������������������������耇�������������������s��6�d�LCKI�8��d�I�STAs�>��_AUTO_DOr��m���IND�D<�δAR_T1�ϿǃT2�������A�X�C� 2(q�cP8�
SONY X�C-56{�u��U��@���� ���А~�H�R5XY ��߭�R5y7����Aff���6�H� $�m��Z� �����������!����E�W�2�{����T{RL�LETE!���T_SCRE�EN �
�kcsc"UD�MMENU 1)�	?  <u�� 1�:o`CLr �������  &_6H�l~ ����/��I/  /2//V/h/�/�/�/ �/�/�/�/3?
??B? {?R?d?�?�?�?�?�? �?�?/OOOeO<ONO �OrO�O�O�O�O�O_ �O_O_&_8_^_�_n_ �_�_�_�_o�_�_o Ko"o4o�oXojo�o�o �o�o�o�o�o5+���_MANUALH߆�DB9�0�����DBG_ERRL�s*���� >����~uqNUMWLIM����dn��ޠDBPXWOR/K 1+���L��^�p������DBT;B_�� ,�}�����u�RqDB_�AWAY}s͡GwCP n�=����_AL
����yr�YGл�n�nx_�p [1-q�́.��
;�y�z�g�����_MM��IS����@A����ONTIM��M�n��ޖ4�
X��I�MOTNEND�M�H�RECORDw 13�� �����G�O�t�b��� ������į֯m�ޯ� t�)���M�_�q��� ���˿:����%� ��Iϸ�m�ܿ�ϣϵ� ��6���Z��~�3�E� W�i��ύ��ϱ� ��� �����z�/��:��� w�������@��� d��+�=�O���s�^�8l�����Oi�������b�M��sN����8���[���)�;�_JX���W����N/�8�9/�k0.:/q/��/���TOLER7ENC��B�>���L��upCSS_�CNSTCY 2�4,���p�/<�� �/??(?>?L?^?p? �?�?�?�?�?�?�? O�O$O6OHO�$DEV�ICE 25�+ І�O�O�O�O�O �O__+_=_O_���#�HNDGD 6��+ՀCzi^LS 27�Ma_�_�_�_�oo'o9oc_�"PA?RAM 8U�%��duKd�$SLAV�E 9�]nW_C�FG :koKcd�MC:\� L�%04d.CSV�Jo<�c�ofr+"A &sCHp�Q��Kn(*_}g�KfOr|q��zyyq�`JP�Ьsk~<�ρ�lRC_OUT ;�M�ρOo_SGN �<K�4��a01�-APR-23 14:35p+�=���F V�t��g�c�Knd���mE�@�S�Þ�ǧj�x�z��cVE�RSION ��V4.0.�1��EFLOGI�C 1=�+ 	�x�`��q���PROG_ENB�)��V2�ULS� ��V�_ACCL{IM���c��q�WRSTJN`ɐ�3��a�MO;��uq�b��INIT c>�*K��a ��wOPT�` ?	��Ȓ
 	R5�75Kc�74!�6"�7"�50F�ׄL��2"��xp�އ��TO�  �z�ů߆V.֐DEX��d���p�ݣPATH A�A\˯*�<���+HCP_CLN�TID ?�c� �{G#|��!I�AG_GRP 2�C�i Q�	 ��ؿÿ��� ��D����mp1m1�0 890123�4567n���=�� ?ϜϮω������r������!�3���\�n����q�G� �߻ߙ�����{���� 9�K�)�o���U�g� ������������3� Y�7�i����+�u��� ������/g yW��9��� 	�-?�>χ :ϫ����|����;/&/_/�˰_O 4Q/�/A/#�/g�/ ?!?혒$-?W?�/g? �?o?�?�?m�?E/O �?ODO/OhOSO�OwO �O�O�O�O�O
_�O._�_R_��<�p c_�_�_C_�_�_�_ �_�_o0o�_@ofoQo��ouo�o�o�o��CT�_CONFIG �D��ʓ]��eg�u��STB_F_TTS��
J��)s��}�xq<v�pM�AU��?�Q�MSW�_CF�`E��  ���OCVIEWfPpF�}�a���� ����*�<���� e�w���������N�� ����+�=�̏a�s� ��������͟\��� �'�9�K�ڟo����� ����ɯX�����#� 5�G�Y��}������� ſ׿f�����1�C�,Uϡ|RC�sG]r!�c΍��ϱ������
���.�tSBL_�FAULT H��ʥxH�GPMSK�2w[��`TDIAG' Iy�qUt���UD1: 6�78901234!5��x��c�P�o�� ��*�<�N�`�r�� ������������;�Vp���@8r��\�>�fTRECP�ߣ�
�ԣ����������� 1CUgy� ������	0��B�?f�UMP_OPTION2pT�a�TR�r3sX��P�ME1uuY_TE�MP  È�g3B�Vp��A��UNInp4u����YN_BRK �J��bEDIT_~y�ENT 1K��?  ,&�R/0P@/}/P�l/�/ �/�/�/�/?�/'?? K?]?D?�?h?�?�?�? �?�?�?�?�?5OOYO @OhO�OvO�O�O�O�O �O_�O1_C_*_g_N_��_r_ MGDI_�STA��q�%N�C�S1L�{ �P�_�_P
Pd7 Yoko}o�o�o�o�o�o �o�o1CUg y������� �� �.�Fa.�T�f� x���������ҏ��� ��,�>�P�b�t��� ������6������ #�=�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ۟���	��5�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�ӿ����� �-�#�I�[�m��� ������������!� 3�E�W�i�{������� ����������7�A Sew����� ��+=Oa s��������� ///9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?��?�?�?O'/1O COUOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�?�_�_ �_oOo;oMo_oqo �o�o�o�o�o�o�o %7I[m� ��_����o)o 3�E�W�i�{������� ÏՏ�����/�A� S�e�w�������џ ����!�+�=�O�a� s���������ͯ߯� ��'�9�K�]�o��� �����ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߷��� ��������-�?�Q� c�u��������� ����)�;�M�_�q� �����ߝ�������	� ��%7I[m� ������! 3EWi{����� ����///A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?���?�?�?�? /O'O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�? �_�_�_�_Ooo1o CoUogoyo�o�o�o�o �o�o�o	-?Q cu��_���� �_��)�;�M�_�q� ��������ˏݏ�� �%�7�I�[�m��� ����ǟٟ���!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ������� ��'�9�K�]�o�� ���߷���������� #�5�G�Y�k�}��� ������������1� C�U�g�y��ߝ����� ������	-?Q cu������ �);M_q ��y������/ /%/7/I/[/m//�/ �/�/�/�/�/�/?!? 3?E?W?i?���?�? �?y?��?OO/OAO SOeOwO�O�O�O�O�O �O�O__+_=_O_a_ {?�?�_�_�_�_�?�_ oo'o9oKo]ooo�o �o�o�o�o�o�o�o #5GYk�_�� ���_����1� C�U�g�y��������� ӏ���	��-�?�Q� c�}���������ɟ ���)�;�M�_�q� ��������˯ݯ�� �%�7�I�[�u�g��� ����ϟ�����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�m���ߛ߭߿�ٿ ������+�=�O�a� s����������� ��'�9�K���w߁� �������������� #5GYk}�� �����1 CUo�y����� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?gU? �?�?�?��?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_�3_E__? �$EN�ETMODE 1�M�5� W o0o0j5��_�[nPRROR_PROG %{Z�%i6�_�Y�UTAB_LE  {[�?�-o?oQo_g�RSEV�_NUM �R  ��Q�`�Q�_AUTO_EN�B  �U�S�T_;NO�a N{[�Q}�b  *��`���`��`��`�`+��`�o�dHIS�}cm1�P�k_ALMw 1O{[ �j4�li0+�� ����_vb�`  {[�a�R2��nPTCP_VER� !{Z!�_�$�EXTLOG_R�EQ3v�i��SsIZ���STK����e�TOL�  m1Dz;r��A �_BWD��瀠f��R��DI�� P�5���Tm1�STEP�)�;�nPU�OP_D�ȌlQFDR_G�RP 1Q{Y�ad� 	-�ʟ�P����E%�ڭ?��#��[���� �
� ��������!��D� /�h�S���w�������@�ѯ
���.��W
$� ]�fvM�����������B�  �A�  @�33��UO��Ϳ��9�$�F�6 F@]��[�g�"σ�F� ?�  �Ϙ�<P����;O��9 �n���r���q�FE�ATURE R��5��QArcTool D��m2Engli�sh Dicti�onaryO�4D� Standar�dH�Analog� I/OG�AZ�e� Shift��r�c EQ Pro�gram Sel�ect��Soft�par����Wel�d��cedureys��@�Core���?�Rampingn��uto��wa'�UpdateM�m�atic Bac�kupM�{�gro�und Edit�E�R�Cameraz��F��Cell�����nrRndIm����ommon �calib UI�����sh�����c�&�.���neC�.�t%y��s����n���Monitorb��ntr>�eliayb��N�DHCPD����ata Acq�uis���iag�nosw����oc�ument Vigewe���ua#��heck Saf�ety	�R�han�� Rob��rvB��qF
�N�ks" �F��(�R�xt w�eavx�chJ�x�t. DIO$�nsfiG� endS Err��L��%s�	r���  �L��FCTN Men�u; �  TP I�nfac(�R�G�en��l�Eq �L�]��p Ma�sk ExcO g�HTJ��xy �Sv#�igh-wSpeS Ski������$�mmuni�cv�on�Hou�r1����Mco�nn}�2(ncr�Lstruc�M�K�AREL Cmd7. L�ua�E#�Run-Ti� E�nv;(_�+z�s�x�S/WO�Lic�ense5"� B�ook(Syst�em)L�MACR�Os,�/Off;se�MMR�����MechStoEp��t�����%i����6xS ��x�1>od��wit�T8�����.$�r;Optm8�?�#��fil"�'�g��%ulti-�T�E�P�PCM 'fun4'�9o��6�E�MRegi� r,��6ri F
KRF���Nu����nH��Adju�hN�Ҵ٦MtatuNA�O
QշRDMUot`�s�covei��Eem0�nw��ERZ� N^ues��9Wo$��_0N�SNPX b�"H�SNJCli}^��urhӝ_z�Q %4ujUo� t1ssagE�jU�A��{_F� U��!n/I|KeMILIB;o~bP Firm^�:%nP1Acc�����TPTX��del�n� XoaA��%&mo�rIP SimulQa����fu� P]��j���3&��ev�.eV�ri3 �o?USB po����iP� a bunexceptS P(DXbu�uVC�r��8V���rvo�u�[��{S�PSC�e
�S�UIK�W� �8<�b Pl�FX�Z�� �M�#�FQ�xuvn�ԇGrid
Qplay΍"`��eR�r.wڊ�RC��g�100iD/1�450��larm Cause/P�edj�Ascii���Load" v�U3pl����yc��k"0Y@Pp@ %RAp��<l�"�NRTL�oS��Online Hel���6L�6L@IA��trG�64MB� DRAM��\�F�ROe���tl!�0.�L�mai#��[�L%�Supmr�1NIР� �cro�LS�U���V�Rmi܉�vrt2SK���O�W� i�������̿ÿտ� ���%�/�\�S�eϒ� �ϛ��Ͽ�������� !�+�X�O�aߎ߅ߗ� �߻���������'� T�K�]������� ���������#�P�G� Y���}����������� ����LCU� y������� H?Q~u� ������// D/;/M/z/q/�/�/�/ �/�/�/�/	??@?7? I?v?m??�?�?�?�? �?�?OO<O3OEOrO iO{O�O�O�O�O�O�O __8_/_A_n_e_w_ �_�_�_�_�_�_�_o 4o+o=ojoaoso�o�o �o�o�o�o�o0' 9f]o���� ����,�#�5�b� Y�k�������Ώŏ׏ ���(��1�^�U�g� ������ʟ��ӟ��� $��-�Z�Q�c����� ��Ư��ϯ�� �� )�V�M�_�������¿ ��˿����%�R� I�[ψ�ϑϾϵ��� ������!�N�E�W� ��{ߍߺ߱������� ���J�A�S��w� ����������� �F�=�O�|�s����� ��������B 9Kxo���� ���>5G tk}����� /�/:/1/C/p/g/ y/�/�/�/�/�/ ?�/ 	?6?-???l?c?u?�? �?�?�?�?�?�?O2O )O;OhO_OqO�O�O�O �O�O�O�O_._%_7_ d_[_m_�_�_�_�_�_ �_�_�_*o!o3o`oWo io�o�o�o�o�o�o�o �o&/\Se� �������"� �+�X�O�a������� �����ߏ���'� T�K�]����������� �۟���#�P�G� Y���}��������ׯ ����L�C�U��� y�������ܿӿ�� 	��H�?�Q�~�uχ� �ϫ���������� D�;�M�z�q߃ߝߧ� ������
���@�7� I�v�m�������� ������<�3�E�r� i�{����������� ��8/Anew ������� 4+=jas�� �����/0/'/ 9/f/]/o/�/�/�/�/ �/�/�/�/,?#?5?b? Y?k?�?�?�?�?�?�? �?�?(OO1O^OUOgO �O�O�O�O�O�O�O�O�$_Q  OH541S?Q2DVoR782EW50EUoJ614iW76EU�AWSPQW1�WRkCRuX8�VTU�V�J545iX�VVC{AMEUCLIO�V�RI�WUIFQV6��WCMSCh�VS�TYLiW2�VCN�REQV52�VR6�3PWSCHEUDO�CVqfCSUEUO{RS�VR869iW�0tW88DVEIO�fR54\VR69��VESET�W�WJ�YWMGEUMAS�KEUPRXY5h7&EVOC�V�`3�X\VX�`hXgX53�fH^xwLCHvOPLv�J50HvPS�wM�C�W�p�g55tVMgDSW�w;wOP;wMPR�Va`0v�`hVPCMg0��`tW�50�51�W51�P�0�VPRS�g6�90vFRD�VRMsCN)f�hH93hV�SNBAg_wSH�LB)fM߇a`XgNuNlx2hVHTC�V�TMI4fYP�fTP�AfTPTX�EL���p�g8[WYPDVwJ95�VTUT<w�950vUECvU�FR�VVCC��O�VVIP4fCSC�L��`I�xtVWEB��VHTT�W6WgW�IO��CG�IG��IPGS=�RC�4fHZXR66�VRU7�gRN�2HvRjz�40vu�tV`DVNV�D�fD0��F�C�TO�WNN0vOL�'hENDQVL×S;LM�fFVRe X K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩπ����������'��  H54�1)�C�2H�R78�2I�50I�J61�4y�76I�AWSuPY�1��RCR���8��TU��J54y5yܘ�VCAMI�oCLIO�RI��UIFY�6��CM�SCY��STYLzy�2��CNREYڻ52��R63X�S{CHI�DOCV��wCSUI�ORS�گR869y�0��8�8H�EIOh�R5�4h�R69��ES�ET�۷�J��WM�GI�MASKI�P�RXY��7I�OC(��3��hڅ�x�w��53�HLCH��OPL��J506��PSgMC��u ���55��MDSW���OP��MPR�(�����%�x�PCMbH�0����50[51��51X0�ڷPRSx�69��F{RD�RMCNy���H93x�SNByAI�SHLBy�M+���NN(2�x�HTC��TMI���e��TPAh�T7PTXi*EL�u ��8g�e�H�J95n��TUT��95��wUEC��UFR��VCC8<O��VI�P��CSC�*��I�i��WEB��HTuT��6��WIO�:�CG�;IG�;IP[GS�:RC��HfܷR66��R7g�R*V2��R&4��5@���U�H�NVDx�Du0�KF�LCTO���NN��OLw�ENuDY�LG;SLMx�FVRh�(�O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o�o�o�o# 5GYk}��� ������1�C� U�g�y���������ӏ ���	��-�?�Q�c� u���������ϟ�� ��)�;�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/�A�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� ������������ �'�9�K�]�o����� ������������# 5GYk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ����������%�1�STD~,�LANGM� H�`�r߄ߖߨߺ��� ������&�8�J�\� n����������� ���"�4�F�X�j�|� �������������� 0BTfx�� �����, >Pbt���� ���//(/:/L/�^$RBTL�OPT�Nu/�/�/�/�/�+DPNK��/�/??/? M�$�S?e?w?�?�?�? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q���������˟ݟ ���%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ����� /�A�S�e�wωϛϭ� ����������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy�� �����	- ?Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O__�99'U�$F�EAT_ADD �?	���TQ~\P  	$X e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������#�5GGTDEMO �RTY   $X������ ��///&/8/R/\/ �/�/�/�/�/�/�/�/ �/+?"?4?N?X?�?|? �?�?�?�?�?�?�?'O O0OJOTO�OxO�O�O �O�O�O�O�O#__,_ F_P_}_t_�_�_�_�_ �_�_�_oo(oBoLo yopo�o�o�o�o�o�o �o$>Hul ~������� � �:�D�q�h�z��� ����ݏԏ��
�� 6�@�m�d�v������� ٟП����2�<� i�`�r�������կ̯ ޯ���.�8�e�\� n�������ѿȿڿ� ���*�4�a�X�jϗ� �Ϡ����������� &�0�]�T�fߓߊߜ� �����������"�,� Y�P�b������� ��������(�U�L� ^��������������� �� $QHZ� ~�������  MDV�z� ������// I/@/R//v/�/�/�/ �/�/�/�/??E?<? N?{?r?�?�?�?�?�? �?�?
OOAO8OJOwO nO�O�O�O�O�O�O�O __=_4_F_s_j_|_ �_�_�_�_�_�_oo 9o0oBooofoxo�o�o �o�o�o�o�o5, >kbt���� ����1�(�:�g� ^�p�������ӏʏ܏ �� �-�$�6�c�Z�l� ������ϟƟ؟��� )� �2�_�V�h����� ��˯¯ԯ���%�� .�[�R�d�������ǿ ��п���!��*�W� N�`ύτϖ��Ϻ��� ������&�S�J�\� �߀ߒ߿߶������� ��"�O�F�X��|� ������������ �K�B�T���x����� ��������G >P}t���� ��C:L yp������ 	/ //?/6/H/u/l/ ~/�/�/�/�/�/?�/ ?;?2?D?q?h?z?�? �?�?�?�?O�?
O7O .O@OmOdOvO�O�O�O �O�O�O�O_3_*_<_ i_`_r_�_�_�_�_�_ �_�_o/o&o8oeo\o no�o�o�o�o�o�o�o �o+"4aXj� �������'� �0�]�T�f������� ��������#��,� Y�P�b����������� ������(�U�L� ^������������ܯ ���$�Q�H�Z��� ~��������ؿ�� � �M�D�Vσ�zό� �ϰ��������
�� I�@�R��v߈ߢ߬� ���������E�<� N�{�r�������� �����A�8�J�w� n������������� ��=4Fsj| ������ 90Bofx�� �����/5/,/ >/k/b/t/�/�/�/�/ �/�/�/?1?(?:?g? ^?p?�?�?�?�?�?�? �? O-O$O6OcOZOlO �O�O�O�O�O�O�O�O )_ _2___V_h_�_�_ �_�_�_�_�_�_%oo .o[oRodo~o�o�o�o �o�o�o�o!*W N`z����� ����&�S�J�\� v����������ڏ����"�O�F�r�  i��������� П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^>p  qk �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |������� ��0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� \�n������������� ����"4FXj |��������0BTfvzm����� ��/ /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo jo|o�o�o�o�o�o�o �o0BTfx �������� �,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx ������� ,>Pbt�� �����//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x���$FEAT_D�EMOIN  V{�����~���_INDEX��������ILECOM�P S����ޑ����ԐS�ETUP2 T�ޕ��  �N �ѓ_AP2�BCK 1Uޙ  �)y�G�V�%=�z�~��h��� {�<�ѯ`������+� ��O�ޯs������8� Ϳ߿n�ϒ�'�9�ȿ ]�쿁�ώϷ�F��� j���ߠ�5���Y�k� �Ϗ�߳���T���x� ���C���g��ߋ� ��,���P������� ��?�Q���u����(� ����^�����)�� M��q��6� �l�%�2[ ���D�h �/�3/�W/i/� �//�/@/�/�/v/? �//?A?�/e?�/�?�? *?�?N?�?�?�?O�?@=O�?JOsO�!�P%�� 2:�*.V1RzO�O2@*�O�O`/C�O_E�@PC_|H_2@FR6:3_"t^_�_'[T���_ �_]U�_�\���_o F�*.F�OOo1A	�_S=o|lo�o/kSTM�o�o\RbP�o }�o$/kH�oW�g�E�0jGIF ���e���-�0jJPG7�a��eM�
����(ZJS���2@�w�ҏ��%
Ja�vaScript�;�CS�h��fU��� %Casc�ading St�yle Shee�ts��@
ARGNAME.DTß
&L�`\ן�������ğ�DISP*���`[���*������H�
TPEIN�S.XML˯w�:�\߯����Cust�om Toolb�ar �O�PASS�WORD��$NF�RS:\c�"� %�Passwor�d Config ���?�|��#�YOG� ֿk�}�ϡ�0����� f��ϊ�߮���U��� y��r߯�>���b��� 	��-��Q�c��߇� ��:�L���p���� ��;���_������$� ��H�����~���7 ����m��� �� V�z!�E� i{
�.�Rd ��/�/S/�w/ /�/�/</�/`/�/? �/+?�/O?�/�/�?? �?8?�?�?n?O�?'O 9O�?]O�?�O�O"O�O FO�OjO|O_�O5_�O ._k_�O�__�_�_T_ �_x_oo�_Co�_go �_o�o,o�oPo�o�o �o�o?Q�ou ��:�^��� )��M��F������ 6�ˏݏl����%�7� Ə[���� ���D� ٟh�ҟ���3�W� i��������ïR�� v������A�Яe��� ^���*���N������ Ϩ�=�O�޿s�ϗ� &�8���\��π���'� ��K���o߁�ߥ�4� ����j��ߎ�#�����Y�;��$FILE�_DGBCK 1�U��F���� < ��)
SUMMAR�Y.DGc��M�D:�����D�iag Summ�ary����
CONSLOG�������[���Console log\����	TPACCN�Q���%������T�P Accoun�tin}���FR�6:IPKDMPO.ZIP�
'�`����Excep�tiond��MEMCHECK���8����o�Mem�ory Data��;�(YF)	FTPN�?�C��q�mment �TBDl;�L =��)ETHERNETa������Ethern�et s�figu�ra���VDCSVRF`FXq/��%6  verify allt/�>�M+�1%DI�FFi/O/a/�/� {%�(diff�/��'�6 CHG01 �/�/�/{?�!?�?�"*f992q?X?j?�?
?�?�?@23�?�?�?��O O�O9F�VTRNDIAG.LS�O`OrO_���A ��nost�ic_>�T6a�)UPDATE�S.MP3_�FR�S:\K_�]��U�pdates L�ist�_�PSRBWLD.CM�_��wR�_�_p�PS�_ROBOWEL����AHADO�W�O�O�O�o�S�hadow Ch�anges�o{qQbNOTI;/�lo~o�Not�ific"�o;�+@AG��j�9� �����w��� B��f�x����+��� ҏa��������'�P� ߏt������9�Ο]� ����(���L�^�� �����5���ܯk� � ��$�6�ůZ��~��� ���C�ؿ�y�ϝ� 2���?�h�����ϰ� ��Q���u�
�߫�@� ��d�v�ߚ�)߾�M� ���߃���<�N��� r����7���[��� ���&���J���W��� ���3�����i����� "4��X��|� �A�e��0 �Tf���� O�s//�>/� b/�o/�/'/�/K/�/ �/�/?�/:?L?�/p? �/�?�?5?�?Y?�?}? �?$O�?HO�?lO~OO �O1O�O�OgO�O�O _ 2_�OV_�Oz_	_�_�_ ?_�_c_�_
o�_.o�_ Rodo�_�oo�o�oMo �oqo�o<�o` �o��%�I�� ��8�J��n�� ��!���ȏW��{�� "���F�Տj�|���� /�ğ֟e�������� +�T��x������=� үa������,���P� b�񯆿���9���� o�ϓ�(�:�ɿ^�� �ϔ�#ϸ�G�����}πߡ�6���C�l�N���$FILE_FR�SPRT  ���V�������MDONL�Y 1U��N�� 
 �)MD�:_VDAEXTP.ZZZs�$����
�6%NO� Back fi�le ��N�S�6�\��߀�Iߍ�� ����i������4��� X�j���������S� ��w���B��f ����+�O�� ��>P�t �'��]��/ (/�L/�p/�//�/�5/�/�/��VISB�CK�؝���*.�VD�/'?� FR�:\� ION\DOATA\?�"� �Vision VD(�S?a/�?�?�/ �?�/�?�?O+O�?OO �?sO�OO�O8O�O\O nO_�O'_9_�O]_�O �__�_�_F_�_j_�_ o�_5o�_Yo�_�_�o o�o�o�o�oxo�o C�og�o��,��P�t��{�L�UI_CONFIoG V��	1>&� $ ��� q���������ˏݏ��$ |x��!�3� E�W�g����������� ҟi����,�>�P� �t���������ίe� ���(�:�L��p� ��������ʿa�� � �$�6�H�߿l�~ϐ� �ϴ���]������ � 2�D���h�zߌߞ߰� ��Y�����
��.��� ?�d�v����C��� ������*���N�`� r�������?������� &��J\n� ��;���� "�FXj|�� 7����//� B/T/f/x/�/!/�/�/ �/�/�/?�/,?>?P? b?t?�??�?�?�?�? �?O�?(O:OLO^OpO �OO�O�O�O�O�O _ �O$_6_H_Z_l_~__ �_�_�_�_�_�_�_ o 2oDoVohozoo�o�o �o�o�o}o�o.@ Rd�o����� �y��*�<�N�`� ���������̏ޏu� ��&�8�J�\�󏀟 ������ȟڟq���� "�4�F�X��|�����в�į֯f��|��$FLUI_DA�TA W��}��j����RESULT �2X�0� �T���L�^�p� ��������ʿܿ� � �$�j�9�L�^�pς� �Ϧϸ������� ���$�6�G�?j�0���~�i�{��r��߱��������� ��/�A�S�e�w�6� �ߡ�������������1�C�U�g�y�j� 
�yߟ�]߿������� 
.@Rdv� ������� *<N`r��� �������/��8/ J/\/n/�/�/�/�/�/ �/�/�/?"?�F?X? j?|?�?�?�?�?�?�? �?OO�?O/cO%/ 'O�O�O�O�O�O�O_ _,_>_P_b_t_3?�_ �_�_�_�_�_oo(o :oLo^opo/O�oSO�o �o�_�o $6H Zl~�����_ ��� �2�D�V�h� z��������o�o�o ���o@�R�d�v��� ������П����� �<�N�`�r������� ��̯ޯ���ӏ� ��A�k�-�������ȿ ڿ����"�4�F�X� j�)��Ϡϲ������� ����0�B�T�f�%� 7�I�[��������� �,�>�P�b�t��� ���{�������(� :�L�^�p��������� ���ߛ߭���6H Zl~����� ����2DVh z������� 
//������a/#�/ �/�/�/�/�/�/?? *?<?N?`?q?�?�? �?�?�?�?OO&O8O JO\OnO-/�OQ/�Ou/ �O�O�O_"_4_F_X_ j_|_�_�_�_�_�O�_ �_oo0oBoTofoxo �o�o�o�oO�o�O �O,>Pbt�� ��������_ :�L�^�p��������� ʏ܏� ���o3��o W��������Ɵ؟ ���� �2�D�V�h� '�������¯ԯ��� 
��.�@�R�d�#��� G����������� *�<�N�`�rτϖϨ� ��y�������&�8� J�\�n߀ߒߤ߶�u� �������Ͽ4�F�X� j�|���������� �����0�B�T�f�x� �������������� �����5_!�� �����( :L^����� ��� //$/6/H/ Z/+=O�/s�/ �/�/? ?2?D?V?h? z?�?�?�?o�?�?�? 
OO.O@OROdOvO�O �O�O�O}/�/�/_�/ *_<_N_`_r_�_�_�_ �_�_�_�_o�?&o8o Jo\ono�o�o�o�o�o �o�o�o�O�O�OU _|������ ���0�B�T�oe� ��������ҏ���� �,�>�P�b�!��E ��iΟ�����(� :�L�^�p��������� ɟܯ� ��$�6�H� Z�l�~�������s�տ ������ �2�D�V�h� zόϞϰ��������� 
�ɯ.�@�R�d�v߈� �߬߾��������ſ '��K������ ����������&�8� J�\�߀��������� ������"4FX �y;��s��� �0BTfx ���m����/ /,/>/P/b/t/�/�/ �/i���/?�(? :?L?^?p?�?�?�?�? �?�?�? O�$O6OHO ZOlO~O�O�O�O�O�O �O�O�/?�/)_S_? z_�_�_�_�_�_�_�_ 
oo.o@oRoOvo�o �o�o�o�o�o�o *<N__1_C_� g_�����&�8� J�\�n�������coȏ ڏ����"�4�F�X� j�|�������q�� ����0�B�T�f�x� ��������ү����� �,�>�P�b�t����� ����ο���ß՟ �I��pςϔϦϸ� ������ ��$�6�H� �Y�~ߐߢߴ����� ����� �2�D�V�� w�9ϛ�]��������� 
��.�@�R�d�v��� ������������ *<N`r��� g�������&8 J\n����� �����"/4/F/X/ j/|/�/�/�/�/�/�/ �/�?�???x? �?�?�?�?�?�?�?O O,O>OPO/tO�O�O �O�O�O�O�O__(_ :_L_?m_/?�_�_gO �_�_�_ oo$o6oHo Zolo~o�o�oaO�o�o �o�o 2DVh z��]_�_�_�� �_�.�@�R�d�v��� ������Џ��o� *�<�N�`�r������� ��̟ޟ���� G�	�n���������ȯ گ����"�4�F�� j�|�������Ŀֿ� ����0�B���%� 7���[���������� �,�>�P�b�t߆ߘ� W�����������(� :�L�^�p����e� wω�����$�6�H� Z�l�~����������� ���� 2DVh z������� ������=��dv� ������// */</��M/r/�/�/�/ �/�/�/�/??&?8? J?	k?-�?Q�?�? �?�?�?O"O4OFOXO jO|O�O�O�?�O�O�O �O__0_B_T_f_x_ �_�_[?�_?�_�?o o,o>oPoboto�o�o �o�o�o�o�o�O( :L^p���� ����_��_3��_ �l�~�������Ə؏ ���� �2�D�h� z�������ԟ��� 
��.�@��a�#��� ��[���Я����� *�<�N�`�r�����U� ��̿޿���&�8� J�\�nπϒ�Q���u� ���ϫ��"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� ���;���b�t����� ����������( :��^p���� ��� $6�� ��+��O���� ��/ /2/D/V/h/ z/�/K�/�/�/�/�/ 
??.?@?R?d?v?�? �?Yk}�?�OO *O<ONO`OrO�O�O�O �O�O�O�/__&_8_ J_\_n_�_�_�_�_�_ �_�_�?�?�?1o�?Xo jo|o�o�o�o�o�o�o �o0�OAfx �������� �,�>��__�!o��Eo ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~���O���s�կ ����� �2�D�V�h� z�������¿Կ濥� 
��.�@�R�d�vψ� �ϬϾ����ϡ��ů '����`�r߄ߖߨ� ����������&�8� ��\�n������� �������"�4���U� �y���O�������� ��0BTfx �I����� ,>Pbt�E� ��i�����//(/ :/L/^/p/�/�/�/�/ �/�/� ??$?6?H? Z?l?~?�?�?�?�?�? ���O/O�VOhO zO�O�O�O�O�O�O�O 
__._�/R_d_v_�_ �_�_�_�_�_�_oo *o�?�?OO�oCO�o �o�o�o�o&8 J\n�?_��� ����"�4�F�X� j�|���Mo_oqoӏ�o ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί௟���Ï%� �L�^�p��������� ʿܿ� ��$��5� Z�l�~ϐϢϴ����� ����� �2��S�� w�9��߰��������� 
��.�@�R�d�v�� �߬���������� *�<�N�`�r���Cߥ� g�������&8 J\n����� ����"4FX j|������� ���/���T/f/x/ �/�/�/�/�/�/�/? ?,?�P?b?t?�?�? �?�?�?�?�?OO(O �IO/mOOC?�O�O �O�O�O __$_6_H_ Z_l_~_=?�_�_�_�_ �_�_o o2oDoVoho zo9O�O]O�o�o�O�o 
.@Rdv� �����_��� *�<�N�`�r������� ��̏�o�o�o��#��o J�\�n���������ȟ ڟ����"��F�X� j�|�������į֯� ����ݏ���u� 7�������ҿ���� �,�>�P�b�t�3��� �ϼ���������(� :�L�^�p߂�A�S�e� �߉��� ��$�6�H� Z�l�~������� ����� �2�D�V�h� z������������ߥ� ����@Rdv� ������ ��)N`r��� ����//&/�� G/	k/-�/�/�/�/ �/�/�/?"?4?F?X? j?|?�/�?�?�?�?�? �?OO0OBOTOfOxO 7/�O[/�O/�O�O_ _,_>_P_b_t_�_�_ �_�_�_�?�_oo(o :oLo^opo�o�o�o�o �o�O�o�O�O�oH Zl~����� ��� ��_D�V�h� z�������ԏ��� 
���o=��oa�s�7� ������П����� *�<�N�`�r�1����� ��̯ޯ���&�8� J�\�n�-�w�Q���ſ ������"�4�F�X� j�|ώϠϲ��σ��� ����0�B�T�f�x� �ߜ߮����ɿ���� �ٿ>�P�b�t��� ������������� :�L�^�p��������� ������ ������ �i+����� �� 2DVh '�������� 
//./@/R/d/v/5 GY�/}�/�/?? *?<?N?`?r?�?�?�? �?y�?�?OO&O8O JO\OnO�O�O�O�O�O �/�/�/_�/4_F_X_ j_|_�_�_�_�_�_�_ �_o�?oBoTofoxo �o�o�o�o�o�o�o �O;�O_!_�� �������(� :�L�^�p�������� ʏ܏� ��$�6�H� Z�l�+��O��s؟ ���� �2�D�V�h� z�������¯����� 
��.�@�R�d�v��� ������}�߿���ş ǿ<�N�`�rτϖϨ� ����������ӯ8� J�\�n߀ߒߤ߶��� �������Ͽ1��U� g�+ߎ��������� ����0�B�T�f�%� �������������� ,>Pb!�k�E� ��{���( :L^p���� w��� //$/6/H/ Z/l/~/�/�/�/s� ��/?�2?D?V?h? z?�?�?�?�?�?�?�? 
O�.O@OROdOvO�O �O�O�O�O�O�O_�/ �/�/�/]_?�_�_�_ �_�_�_�_oo&o8o Jo\oO�o�o�o�o�o �o�o�o"4FX j)_;_M_�q_�� ���0�B�T�f�x� ������moҏ���� �,�>�P�b�t����� ����{����(� :�L�^�p��������� ʯܯ� ����6�H� Z�l�~�������ƿؿ ����͟/��S�� zόϞϰ��������� 
��.�@�R�d�uψ� �߬߾��������� *�<�N�`�ρ�Cϥ� g���������&�8� J�\�n���������u� ������"4FX j|���q���� ���0BTfx �������/ ��,/>/P/b/t/�/�/ �/�/�/�/�/?�%? �I?[?/�?�?�?�? �?�?�? OO$O6OHO ZO/~O�O�O�O�O�O �O�O_ _2_D_V_? _?9?�_�_o?�_�_�_ 
oo.o@oRodovo�o �o�okO�o�o�o *<N`r��� g_�_�_���_&�8� J�\�n���������ȏ ڏ����o"�4�F�X� j�|�������ğ֟� ������Q��x� ��������ү���� �,�>�P��t����� ����ο����(� :�L�^��/�A���e� ������ ��$�6�H� Z�l�~ߐߢ�a����� ����� �2�D�V�h� z����oρϓ��� ���.�@�R�d�v��� �������������� *<N`r��� ������#�� G	�n����� ���/"/4/F/X/ i|/�/�/�/�/�/�/ �/??0?B?T?u? 7�?[�?�?�?�?O O,O>OPObOtO�O�O �Oi/�O�O�O__(_ :_L_^_p_�_�_�_e? �_�?�_�?�_$o6oHo Zolo~o�o�o�o�o�o �o�o�O 2DVh z������� �_��_=�O�v��� ������Џ���� *�<�N�r������� ��̟ޟ���&�8� J�	�S�-�w���c�ȯ گ����"�4�F�X� j�|�����_�Ŀֿ� ����0�B�T�f�x� �Ϝ�[�������ϵ� �,�>�P�b�t߆ߘ� �߼������߱��(� :�L�^�p����� ������Ͽ�����E� �l�~����������� ���� 2D�h z������� 
.@R�#�5� �Y�����// */</N/`/r/�/�/U �/�/�/�/??&?8? J?\?n?�?�?�?cu ��?�O"O4OFOXO jO|O�O�O�O�O�O�O �/�O_0_B_T_f_x_ �_�_�_�_�_�_�_�? o�?;o�?boto�o�o �o�o�o�o�o( :L]op���� ��� ��$�6�H� oi�+o��Oo��Ə؏ ���� �2�D�V�h� z�����]ԟ��� 
��.�@�R�d�v��� ��Y���}�߯����� *�<�N�`�r������� ��̿޿𿯟�&�8� J�\�nπϒϤ϶��� ���ϫ��ϯ1�C�� j�|ߎߠ߲������� ����0�B��f�x� ������������� �,�>���G�!�k��� W߼�������( :L^p��S� ��� $6H Zl~�O���s�� ���/ /2/D/V/h/ z/�/�/�/�/�/�/� 
??.?@?R?d?v?�? �?�?�?�?�?��� �9O�`OrO�O�O�O �O�O�O�O__&_8_ �/\_n_�_�_�_�_�_ �_�_�_o"o4oFoO O)O�oMO�o�o�o�o �o0BTfx �I_������ �,�>�P�b�t����� Woio{oݏ�o��(� :�L�^�p��������� ʟܟ���$�6�H� Z�l�~�������Ưد ꯩ��͏/��V�h� z�������¿Կ��� 
��.�@�Q�d�vψ� �ϬϾ��������� *�<���]����C��� ����������&�8� J�\�n���Q϶��� �������"�4�F�X� j�|���M߯�q����� ��0BTfx �������� ,>Pbt�� ������/��%/ 7/�^/p/�/�/�/�/ �/�/�/ ??$?6?� Z?l?~?�?�?�?�?�? �?�?O O2O�;// _O�OK/�O�O�O�O�O 
__._@_R_d_v_�_ G?�_�_�_�_�_oo *o<oNo`oro�oCO�O gO�o�o�O&8 J\n����� ��_��"�4�F�X� j�|�������ď֏�o �o�o�o-��oT�f�x� ��������ҟ���� �,��P�b�t����� ����ί����(� :������A����� ʿܿ� ��$�6�H� Z�l�~�=��ϴ����� ����� �2�D�V�h� zߌ�K�]�o��ߓ��� 
��.�@�R�d�v�� ����������� *�<�N�`�r������� ������������#�� J\n����� ���"4EX j|������ �//0/��Q/u/ 7�/�/�/�/�/�/? ?,?>?P?b?t?�?E �?�?�?�?�?OO(O :OLO^OpO�OA/�Oe/ �O�/�O __$_6_H_ Z_l_~_�_�_�_�_�_ �?�_o o2oDoVoho zo�o�o�o�o�o�O�o �O+�_Rdv� �������� *��_N�`�r������� ��̏ޏ����&��o /	S�}�?����ȟ ڟ����"�4�F�X� j�|�;�����į֯� ����0�B�T�f�x� 7���[���Ͽ����� �,�>�P�b�tφϘ� �ϼ��ύ�����(� :�L�^�p߂ߔߦ߸� �߉�������!��H� Z�l�~�������� ����� ���D�V�h� z��������������� 
.�����s5� ������ *<N`r1��� ����//&/8/ J/\/n/�/?Qc�/ ��/�/?"?4?F?X? j?|?�?�?�?�?��? �?OO0OBOTOfOxO �O�O�O�O�O�/�O�/�_%Y�$FMR2_GRP 1Y%U�� �C4  B��0	 �0c_u\`PF�6 F@�S��Q�T�J`S�_�]`P?�  �_�_<P��a;O��9 n�e�]A`+o=kBH]SB�YPX`;aO@�33ce�\�_<�o�Y@UO߯a�o �_�o�o�o�o4 XC|g����}�9R_CFG ZF[T ��(�|:��{NO FZ/
F0p� u��|�RM_CHKTYP  6Q�0NPPP�P8QROM��_MsIN���3����u�|`X9PSSB�s�[%U aV��5�
���u�TP_DEF_O/W  �4NS1��IRCOM��B���$GENOVRD�_DO���1o�T[HR�� d��du�o_ENBa� u��RAVC?S\Ӈހ ��U"����1��?�P�sj ��ՑOUBPbF\�x�sXF�sU<�� �]ǯq���ᯬ��3C�YP�YP�0%��d��1A@M�?��U�vY��#�֐SM�T?Sc�RP��4���$HOSTC�r1�dFY߀��? 5	
�
�
��6:��9eVχϙ� �Ͻ���u��� ��$��G�H���	anonymousK�yߋ��߯��� 	��-�
� A�c���R�d�v���� ����������M�_� <�N�`�r��������� ����7�&8J \�������� !�3�"4FX�� ��������� //e//T/f/x/�/ ��/��/�/�/?? as���/s?��? �?�?�?�?9/O(O:O LO^O�?�/�/�O�O�O �O�O5?G?Y?_mOZ_ �?~_�_�_�_�_q_�_ �_o oC_Do�Ohozo �o�o�o�O	__-_
 Aoc_@Rdv��_ �����Mo_o <�N�`�r����o�o�o ���7�&�8�J� \����������ُǟ !����"�4�F���챿ENT 1e��� P!ڟ��  ����ï��篪�� ί/��;��d���L� ��p�ѿ�������ܿ �O��s�6ϗ�Zϻ� ~ϐ��ϴ����9��� ]� �Vߓ߂߷�z��� ���������4�Y�� }�@��d����������C��g�*�?QUICC0t�P�b�����1�������2��c!?ROUTERd@�R�!PCJO�G��!19�2.168.0.�10����CAMP�RT�!�1� +RT}/A��h�NAME �!u�!ROBO��S_CFG �1du� ��Auto-s�tarted��FTP��;!͏ϟ f/��/�/�/�/�/o� �/??,?O/=?�/t? �?�?�?�?��/&/8/ OL?n/,O]OoO�O�O Z?�O�O�O�O�O"O�O 5_G_Y_k_}_�_���� ��ʏ_�_BOo1oCo Uogo._�o�o�o�o�o �_xo	-?Qc �_�_�_��o�o� ��)��oM�_�q��� ���:���ݏ��� %�l~������� ��ǟٟ���ď!�3� E�W�i��������ï կ���@�R�d�A�x� e�������������|� ����+�N�O��s� �ϗϩϻ���&�8� :��n�K�]�o߁ߓ� ZϷ���������"ߤ� 5�G�Y�k�}������ �Ϩ����B��1�C� U�g�.���������� ��x�	-?Q���_ERR f��aqPDUSI�Z  ��^����>�WRD �?%���  �guest ����);��SCD_GROUoP 3g, !��� �LOuA��RES��TM� $�T�_�ENBs TT�P_AUTH 1�h� <!i?PendanGR.���A!KAREL:*R/[/m-�KC�/�/�/z �VISION SCETk?�/F!? ?1?w#U?C?m?g?�?��?�?�?�?�>!$CT_RL i�;H���
��FFF�9E3�?��FR�S:DEFAUL�T`LFANU�C Web Server`JNB!$� �	L�O�O�O__,_�oWR_CONF�IG jp��`OqIDL_CPU_PC@���B����P BH�UMIN�\x�U?GNR_IOz������PNPT_S_IM_DO�V�[�STAL_SCR�N�V �6F�QTPMODNTOLg�[�ARTY�X�Q�V�� %  gx�SO�LNK 1k� }�o�o�o�o�o ��bMASTE�P�zi�UOSLAVE� l�AuRAM�CACHE0(bO>'!O_CFGr�cƊsUO0��rCY�CLq�uy@_AS�G 1maW�
 �)�;�M�_�q� ��������ˏݏ��\{�rNUM��	�
�rIPo�wRTRY_CN@�R�
<�ra_UPD��a��� �r�p�rn�P~u��u�PSDT�_ISOLC  �P{v"�J23�_DSrd.N�O�Gg1oP{<���d<�P� ?���R��?��館Q ��̯ޯ𯯯�&�8�J�������*��P�q4i��PhpECso�U�KANJI_*pK��_³� MON pp;_��y�(�:�@L�^�pϒ~"��qa\�EF�ŭ���CL_�L�P'�J�İEYL_OGGIN�pu��F���$LA�NGUAGE ,�FabyD <�q�LG�qr�y�aW ���xu �e�i���P���'0������;��cMCH �;��
��(U�T1:\����  ���������!�3�E�\�i�{��(���l�LN_DISP �sP�ئ�����O�C4b�RDz�S�A�@�OGBOOK tM�d��>A���k�X�܏����������<O�Y���	>F	Q������N`���O�_BUFF [1u�me2kE �j�FB�iG�� G>P}t� �����///�C/��~DCS yw�{�=��� G��/�/�/�/Z$�IO 1x�{ ğ3D��?*?<? N?b?r?�?�?�?�?�? �?�?OO&O:OJO\O�nO�O�O�O�O�O�%E�PTM�dh�#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo�goyo�o-��BSEVt�����FTYP➁_�o�m��R�Sh���|��FL 32y=����/��������(T�P����b'�NG�NAM�6%.�V$UPS��GIh������f�_LOADP�ROG %��%�REQMENU���MAXUAL�RM'��A5�̀l�_PRh��� E�	ˀC��zM��������,�P 2{�� ت	�aڀ	�|�f4��~����� �����(Ο���3�� (�i�T���x���ï�� �ү�� �A�,�e� P�����~������ƿ ؿ��=�(�a�s�V� �ςϻϞϰ������  �9�K�.�o�Zߓ�v� ���ߴ������#�� G�2�k�N�`����� ���������
�C�&� 8�y�d����������������ćDBGDEF |$�:!"��$6 _LDXDI�SAQ�#��#MEM�O_APK�E ?=$�
 H ������"~ˀISC 1}$�%��oy�M�����QE_M?STR ~�m%�SCD 1�� �T/�x/c/�/�/�/ �/�/�/�/??>?)? b?M?r?�?�?�?�?�? �?O�?(OO%O^OIO �OmO�O�O�O�O�O _ �O$__H_3_l_W_�_ {_�_�_�_�_�_o�_ 2ooBohoSo�owo�o �o�o�o�o�o�o. R=va���� �����<�'�`���MJPTCFG 1�+]�%������MIR 1��%Ԁp�@T��q���T�< G ?��%��t �7�q��i������� ������1�C�֟�� j�L�V�x���P����� ί��0�T�E �q� ���8���������� ������ �B�p�R� �ϵ���Z�|���п�� ��6���>�l�R�d߆� �ߖ����ߌߞ���2� ��@�z�`���� ��������+�=����� ���X�b�t������� ������*��o� 6�������� �
@nP� ��Xz���� 4/�,/j/P/b/�/�/����K����� � �/��LTARkM_�"�̅� ��"����6?>4��ME�TPU  T���%��NDSP?_ADCOLX5� �c>CMNTy? ~l5MST ��-��?���!�?�4l5PO�SCF�7�>PR�PM�?�9STw01����4܁<#�
 gA[�gEwO�GcO�O�O �O�O�O�O_�O_G_ )_;_}___q_�_�_�_��_�Ql1SING_�CHK  |?$_MODAQ3�����,�.#eDEV �	��	MC:>WlHSIZEX0�-��#eTASK �%��%$1234?56789 �o�e�!gTRI����� l̅%&�0O2}���cYP�a���9d"cEM_IN�F 1�7;a�`)AT&FVg0E0X�})�q�E0V1&A3&�B1&D2&S0�&C1S0=�})�ATZ�#�
�H@'�O��qCw��A�@��b�ˏ���� � &�������3��� ۏȟڟ������"�4� �X�����A�S�e� ֯៛��C�0���� f�!���q�����s�� ������ͯ>��bϙ� sϘ�K���w������� �ɿۿL����#ϔ� ��Y�����ߩ߳�$� ��H�/�l�~�1ߢ�U� g�yߋ���� �2�i� V�	�z�5����������PoNITOR�0G� ?kk   	?EXEC1�2U2345T�`789���(� 4�@�L�X�@d�p�|�2�U2�2�2�2�U2�2�2�2�U2�3�3�3(�#aR_GRP_S�V 1��{ (`�Q���#a�a_Ds���n�ION_DB�-`�1m�1  ���0qFh"%p0&1��2Gg��N Bl"%}"Fi-ud1}e�/�/�/1PL_N�AME !�e�� �!Defa�ult Pers�onality �(from FD�)b"P0RR2� �1�L68L�@P�!K`
 d �:?L?^?p?�?�?�? �?�?�?�? OO$O6O�HOZOlO~O�O�Oc(2 )?�O�O�O__,_>_P_b_t_f"<�O�_�_ �_�_�_�_
oo.o@o�Rodotl�"Q �_�m
�o�of$P�o�o  $6HZl~�� ������o�o2� D�V�h�z������� ԏ���
��.�@�� !�v���������П� ����*�<�N�`�r�Ą���e����(ïխf"d��� �(�6������y�d���P� ������ Ŀֿ�����:ϐ��h]�m�f"��	`���ϲ��σ�:�o�Ab)�����c' A�  /�	23��)X ����E ���X, @D� M t�?�z�n�?f <|�f!AI�t�jު�;�	l��	 �� � ?�h�Y Z ����� � x � � ������K_K �}K7X�K���J��?J�+�Ƀ�%��ԯC@�6@�
�\��(E@�Sє���.��=�N��������T;f��a������$��*  ´ [ �@ �>����!�z�w�����<�
�����Z!/������yD�  �  �  �`��#  �l����-�	�'� � ���I� �  y�0�&�:�È��?È=�����x�@����%�f���f�(�2�+�a!v�  '�Y��@�!�p@���@j��@��@��C��{C� �� C���C��C��R!��A���=����%"T�Bb $/��Lf!Dz��o��~�@�����R!��A �л�D�  X ,>f �?�ffG�*/</� }�q/�+��8~`�/�*>��H$��(�(~`�%P�(�������>�$�����<�	<S��;�9<���<#*o<���M,@�K;|���f��",�?fff�? ?&�0T�@��.�2�J<?N\��55	��1��(� |��?z��?j7��[/0O OTO?OxOcO�O�O�O`�O�O�O{h�5F�� �O2_�OV_�?w_�9I_ �_E_�_�_�_�_oo oLo7opo[o�oo�o �oU�o�o��m_3�_�Z�o~���O*��& Q/�wl��q
��m.��+�d�V���Aa0��5uCP���L�<č?�����#��Y�/Ӄj6�B]�D��CC3�� z���������@I��l����A���A��PA ��R?�1>��-8��������O\����Q����#�
؞���A�иRA���C;���Q섟�"\)C0����qBo
=���Q�����8�Hp��G�� H�0�H��E1� C�&��Hy��I���H��%F�� �E,�s�]�i�E�I��@H����H��E# D�7�د�կ� ��2��V�A�z�e�w� ����Կ������� @�R�=�v�aϚυϾ� ����������<�'� `�K߄�oߨߺߥ��� �����&��J�5�G� ��k���������� �"��F�1�j�U��� y������������� 0T?x�u� �����tP�(<3�(���	4���<�̷�t�Ӂ3���8����ʭ���Ӂ� &n�
/4�f4yϱ$- $)d/R/�/v/�/�,Յ%PD2P�.�a�o?@Z?=?(?a?L<?g?�n?�?�?�?�?�?  �����?�?+OO OO:OsO?�o�O�O�O�L7�O�O_�O _F_4_JQ�L_^_�_�_p�_�_�_�Z  2jO�o  B��}���Cq���Ӏ@��Rodo@vo�o�o�o�mۃo��o�o/AӄJhDӀӀ�aӀ؎
 I�� ������)�;��M�_�q����sq ����1��"�$�MSKCFMAP�  $%� �Vsqoq莼��ONREL  ��%Ӂ�P��EX_CFENB�
у����FNy�'��JOGOVLIM��d��d��KEY��q�z�_PA�N�������RUN�a���SFSPD�TY� '����SI�GN��T1MO�Tc����_CE_GRP 1�$%Ӄ\dOh�\O�� ���T��ɯ����� #�گG���<�}�4��� ��j�׿�����Ŀ1� �*�g�ϋϝτ��πx���������f��Q?Z_EDIT�͇���TCOM_CF/G 1�ɍ~vv��ߚ�
V�_ARC�_"��%P�T_M�N_MODE���0�UAP_CP�L��4�NOCHE�CK ?ɋ �%�3�E�W�i� {���������������/�A��NO_?WAIT_L�K�66�NT^��ɋu|ޓ�_ERR@�2�ɉ�Q� ���������4F��MO����|ߍ�59<���?����np���PARAuM��ɋ�rv`�3u7�_^ =�P�345678901x��s��� �//�9/K/'+t7��}/�,"�/��ODRDSP���0��OFFSET_C�ARA���&DIS��/�#S_A��AR�K�L�OPEN_FILE0h���L����OPTION_�IO����m0M_P�RG %Ɋ%$�*�?�>I3WO50-�F�0� �5D���2��0@�'A	 ���C���#��� RG_DS�BL  Ʌ��v|rO�!RIENTkTO��!C�mp�ҁ,a� UT_SIM_Du7Ђ��� �V� LCT � ��H��4���I�%y��A�_PEX��?TR[AT�� d0�T>� UP ��N�pK��i_{_XrfS`�bgq�Rn�}]�$��2?��L68L�@P�C
 d�/�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\��2�_������ �
��.��{X�j� |�������ď֏�������� G�X��PX�~��"Pk�����̟ ޟ���&�8�J�\� n�������������� ���"�4�F�X�j�|� ������Ŀֿ���ɯ ۯ0�B�T�f�xϊϜ� ������������,�0>���|�}ߏ�S�$�߿ޤ����׀b�bݢ/3��W�
� @L�v�l�~���� ����J��Q�'�)L�	``�Z�l�~���:�o�A��������>K�A�  ���T��POOP1�[_�v��TH���E=D�X, @D�C  2��,?��D4429�h;��	l�	@� �� �h��� ��� � x � �� ��J�H��H2�-HL���H�lH�WG���=�3Ho��,J�C��@p�@Eז@�P1w#��0�@�S �>P�P%ICUB��< ��K��@��a��y�  ��  �  � #�0�*&�H/��	'� � �f"I� � � ����=��q͊/�+�@�/@� �>A�/M+>B����N�@4?  '�x0L4�0C�@C�W� CC�C��Y?k?D�  ��A�!����������B�@�1�����!
ENz�-O�QO<OaO��O^/p(�1�E�S� ú<��1�P.   �?�ff��O�O��O 7�/_A[sA8��W_eZ>�' I�FjJ(��UP�X��I����#�T[���<�	<S��;�9<���<#*o<���5�\@�	k:���#�R��?fff�?� ?&D`oD@��.Vb�J<?N\�be:��2?aKjI :�o8�o(g~_�o �o�o6!ZE~ �{������ �o�o�o�h����w� ����ԏ��я
���.� �R�=�v�a�?��o� e+��O����<�N�`�r�Z���@_��l� /�ȯ+��ׯ�"����A`>��?��C�s�
�П��?Ƀء����̿n	ĭ/X���B�DF90CC�ޚ��������^�@I�*�����A��A���PA �R?��1>�-�������ÍO\������Q���#�
������AиRA����C;����Q�B��0\)�C0���q�Bo
=��Q�������Hp���G� H�0��H��E1�� C���Hy���I��H��%F�� E,�1���i�EI��@�H���H��E# D��� �ߨߓ��߷������ ��8�#�5�n�Y��}� ������������4� �X�C�|�g������� ��������	B- fxc����� ��>)bM �q�����/ �(//L/7/p/[/m/ �/�/�/�/�/�/?�/ 6?H?3?l?W?�?{?�?@�?�?�?�?O��(��g3�([��T��BE�5�̷�2ODOX��3���^OpO~B��ʭ�O�OX�� &�n�O�O4�f4yϱ�M�I"__F_P4_j_X\��PbP�^�����_O�_�_�_o
l?%o,oeoPouo��o�o  ���� �o�o�o�o�o1�_ ��dR�v|7����������� 
��R�@�v�d������  2(я  B(G�;�G�C/�D�X�@K��"�4�F�X�j�{���������ɟ۟����X���X��X���X���
 �W�i�{������� ïկ�����/�A����1� ���K1���"�$PARA�M_MENU ?��E� � MNU�TOOLNUM[[1]݆��F~������AWEP�CR��.$INC�H_RATE���SHELL_CF�G.$JOB_B�AS߰ WV�WPR.$CEN?TER_RI�������AZIMUTH_ OPTB�����ELEVATIO�N TC����D�W�TYPE S�N�ARCLIN�K_AT �STA�TUSǳ]�__V�ALU߱̰LE}P��.$WP_�� ���U�̢ϴ������� ���7�2�D�V��z��SSREL_ID�  �E�Q���U�SE_PROG �%��%{��ߏ�C�CRT�ԶQ����_HOST !��#!��5���T�P�߈Q��*�S����_?TIMEOU�Ս��  z�GDEB�UG�Љ���GINP_FLMSK��f��TR����PGd��  ����$�CHP����Q���z� tߪ��������� (:c^p��� ���� ;6 HZ�~���� ��// /2/[/��WORD ?	��
 	RS��CPNn�BM3AIW��#SU&��#�TEt�CSTY9L COL0eW(��/W�TRACEC�TL 1��EN�� �P�P7_DT Q��ED0~!0D � �So��QQ6�[;q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k��}�6LEW���5���3  �6_U�P �<;b������ ���&�0��M$a��R�\0R��  ��)_DEFSPD ���{2��  �z��INؐTRL ɡ��a�8!�h�PE�_CONFIܐ�N7���M!b,WLIDٓ���	Ĩ�GRP 1�9� lM!A>f�f��\�
�=D�  DZ�� D
�@�
�M d!�?�O��������H�"�$�i� ������m�B��̱��������̿��&�B34�$�]�o�>Y� <<j��t� ��pϪ�������όπ�O��_߅�p��z�ӳ�M 
���ߊ��� ���5� �Y�D�}�h� ��������������*�)<�
V7.10beta1�� A�k�\��B
��(�Y�?&{ffp�>.{X�
�����X�B�!념�A{33#A�&�(�h� -���P��������pM"��3EWM$ғ��KNOW_M  �0��ȤSV ]�:�%�� �����I�M"G��M�=��(�	������.�* ��7��M#�)�Y�@)���M % .ѐȡMR�=�$�`���f/x+��ST�1 1�<9^ 4�()�o��/�/�/ 
?�/?!?S?E?W?�? {?�?�?�?�?O�?�? >OO/OtOSOeOwO�'�2�,��/���<�O�O� 3�O�O�O�O��'4_-_?_Q_�'5 n_�_�_�_�'6�_�_�_�_�'7o&o8oJo��'8goyo�o�o�'M�AD�� ȕ�EO�VLD  ����P}�$PARNUM  �+?Q�#�SCHy ȕ
�wlq�y��uUPD�l=u���E_CM�P_u����_�'�ݥ%�ER_CHK�3�ۣ �G�0�B�RqSA �ȡ_MOp䕏��_���E_REWS_G� ���
�� p�"��F�9�j�]�o� ����ğ���۟����o��@���1�� PN�m�r��mP���� ����P̯���` �*�/��f`J�i�n��惹`�������V �1���ށ�@]�s8��THR_ICNRA �q]مd�oMASS)� Z=��MN(�[�MON_�QUEUE �P�����!ބN*��Un�NkƔȫ�ENqD��Ώ��EXE�ό���pBE���ϫ�O�PTIO��׋��P�ROGRAM %��%��習��?TASK_It �OCFG ���x��ߵ�DATAx-����G2�$� 6�H�Z�l����� �������� �2��߯INFOx�� ��������������� ��	-?Qcu �������N�Z��� ����pK_�����z�5�G��2�D X�,		x�=�{���@���$a�����0�_EDIT �������WERF�L��Ó#RGADoJ ��AЛ@R$?�]%0�5&��?�����?����A<��z�%��o�/)(/s#2��'"	H��l�|!?8�Aٴw�t$26*A0=/C2 **:L2�??Q3m=���2�5��+1�9��/�? y=�=�?�?�?�?�?KO �?O5O+O=O�OaOsO �O�O�O#_�O�O__ _�_9_K_y_o_�_�_ �_�_�_�_�_goo#o QoGoYo�o}o�o�o�o �o?�o�o)1� Ug������ ��	���-�?�m�c� u����ُϏ�[� ��E�;�M�ǟq��� ������3�ݟ��� %���I�[�������@��ǯ������	�� ��𰄿����39߿53���ϧ�0�B�o'PR�EF �*0�0
5%IORIT�Y:���9!MPD�SP8�'*�"��UT���34&ODUCT����E��&OG_TG$ ������TOENT 1��� (!AF_INE��Y�J�?!tcpdߌݟ!ud{ߴ�!icm���.��kXYx#���1�)� Y1�*�0��S�6�B��f�� �����������!�3� �W�>�{���*��x#��)�"�/�������Y7/c<��44���(�.A�",  �u�(}���+%�^Ŀf�x�,9!�PORT_NUM���0�9!_CARTREP% |�aSKSTA�ǻ 4LGSV������#0Unothing�����L�]TEM�P ����T���_a_seiban�,/�</b/M/ �/q/�/�/�/�/�/�/ �/(??L?7?p?[?�? ?�?�?�?�?�?O�? 6O!OZOEOWO�O{O�O �O�O�O�O�O_2__ V_A_z_e_�_�_�_�_�_�_�_o�VER�SI����M` �disable�d'oSAVE ����	2670/H782J�o�o�!$�o�o���o 	�x��V��.�e@Kt���J�c|��o���mb_� 1����`*�p�!��4�F��W�URGE_ENBЪ�(���WFr�DO���+��WRГ���WRU�P_DELAY ��,��R_HOT %{���#����R_NORMA�L����W�&�SE�MI6�\���U�QS�KIP���#�x o��	o��(��� Y�G�}�����g�ů�� կ�����C�1�g� y���Q���������� 	�Ͽ-��=�c�uχ� Mϫϙ������Ϲ���)��M�_�q����$�RBTIF��0R�CVTMOUEv����DCR�}Ǿ� ����C04^@�����3��띭3����*vJ���-�7���I�4�<��	<S�;��9<��<#*o<��M�Q 7���y���� ����/�A�S�e�w�������RDIO_TYPE  �����EFPOS1W 1�ui� x A
-���G2k�o� *�N���� 1�UgN� ��n��/�/ Q/�u//�/4/�/�/ j/|/�/??;?�/_? �/�??�?�?T?�?x? O�?%O7O�?�?OO�jO�O��OS2 1�ԋZO�O_�Ox6_�O��3 1��O��O�O,_�_�_�_L_S4 1�c_u_�_�_�?o*oco�_S5 1��_
ooVo�o�o�o>voS6 1͍o�o��o�oiT�S7 1�"4F����"��S8 1� ������~���5��SMASK 1����  �� �ՇXN�O���:�D���M�OTE��=�Z�_?CFG �a����A���PL_RAN�G]��ߛ�OWER� �%�ΐ��S�M_DRYPRG %%�%^��ԕTART �ƞ��UME_PRO����p�=�_EXE�C_ENB  <���GSPDI���8���Ѣ�TDB�����RMϯ��IA_O�PTION����\��U�MT_݀T��d_���*�z��9���C�ˀ���𥿷����OBOT�_ISOLC"������ֵNAME� %�_���O�B_ORD_NU�M ?Ƙ���H782  ˄h�@h�$�h����h�>�PC_TI�ME�ם�x��S2�32z�1����L�TEACH ?PENDAN��v��A�~�]�H@M�aintenance Cons˂���ˆ"�DDNo Use~�E�߀i�{ߍߟ߱ߵ���N�PO#���A�!����CH_LL���U���	3���!OUD1:Y� �R܀�VAILI���|��U�SR  %������R_I�NTVAL��������V_DA�TA_GRP 2��%���X�D��P ��W���{�f�%����� ����������$ &8n\���� ����4"X F|j����� ��//B/0/R/x/ f/�/�/�/�/�/�/�/ �/?>?,?b?P?�?t? �?�?�?�?�?O�?(O OLO:O\O^OpO�O�O �O�O�O�O_ _"_H_�6_l_U��$SAF�_DO_PULS���V���X��Q�PCA�N������SC���(�����ˀq����x�C�C�
�˂ p�o0oBo Tofoxoo�o�o�o�oX�o�o�����bHe�!r �dt:ql�(s�� @��fx���~Ny� D�t��_ @�T�������T D��*�S�e�w� ��������я���� �+�=�O�a�s�����^`u2����ǟі��C���;��o2���p����
�t��Di����aC��  � ���Cђax��Qa�s� ��������ͯ߯�� �'�9�K�]�o����� ����ɿۿ����#� 5�G�Y�k�}Ϗϡϳ� ����������1�2��aZ�l�~ߐߢߴ� ������9�u�(�:� L�^�p��������2�0�D��N�	� �-�?�Q�c�u����� ����������) ;M_q���� ���%7I [m����� D��/!/3/E/W/i/ {/�/�/
��/�/�/�/ ??/?A?S?������ r�?�?�?�?�?�?�? O#O5OGOYOgIzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<oNo`o5�艟9�ko�o �o�o�o�o&8 J\n������pj�o��2����S����	12345678+��h!B!�)��4���`��|� ������ď֏���� ��o5�G�Y�k�}��� ����şן����� 1�C�U�f�$������� ��ѯ�����+�=� O�a�s�������h�z� ߿���'�9�K�]� oρϓϥϷ������� �Ͼ�#�5�G�Y�k�}� �ߡ߳���������� �1�C�U��y��� ����������	��-� ?�Q�c�u�������j� ������);M _q������ ���%7I[m ������� /!/3/E/W/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?�?�?�?"�sm��?�?q/O�O*OF�Cz  �Bpqj   ��h2�bm�} �ph
�G�  	��r2�?�O�O�O�O�ok>�_Dlo�<� �OB_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o'_�o�o �o�o(:L^ p�������  ��$�>ISB�1�A�iB<S��$SC�R_GRP 1���8� � �� �SA� dE	 /������� ���1B���SG��ۏɏ��:M�s@��D^@D/^��E��� \�ARC Ma�te 100iD�/1450ҁA�M�ҁMD45� 678SC
1/2345��9��ӅAE����KyBד_�� SF�߃� S��Ó��Ӂ�	yJ6�H�Z�l��~�SD��H���������Əǯ ���Ά�oSAگC�`֯g�N���v�B�M@!Ʋ���ɴ��A^@ؿ�  @S@𵬁@���� ?PŬ�H�M@)�ۺ��F@ F�`S�[�~��j� �ώϳ���������!� ��� �L�7�I�[�m�B�{���߬����� 	����?�*�c�N�� r��_��)������dG�@��0�SB�@P6��6�J���h�p�M@Ȇ��� ��߃�?��SDA���H������ Qƒ�SA 3E��!pht�U (� ������ ��$SF_�EL_DE�FAULT  ~���S@�@HOTSTR�L��`MIPOWERFL  BExX?�WFDOM� �RVENT? 1�����w� L!DUM�_EIP.���j�!AF_INExL/SD!FT��@./d/!���/ ��S/�/!RP?C_MAIN�/�(q��/�/�#VIS�/�)��/H?!TP&;0PU??�d7?�?�!
PMON_POROXY�?�e�?��?[2�?�f�?,O!�RDM_SRV�-O�gOxO!RȲ��O�hgO�O!
�� M�?�i�O_!RLSYNC_���8�O\_!R3OS��\�4K_�_�!
CE]0MTC�OM�_�k�_�_!=	�RCONS�_��l�_@o!�RWA'SRCGO�m/o�o;!�RUSB�o�n{o�ow/�o;C�o�o %Jn5�Y��:RVICE_K�L ?%� (�%SVCPRG1����u2�
��p3-�2��p4U�Z��p5}����p6�����p�7͏ҏ�p����9�"��t�OJ��q� r��q����qG��q o���q����q��:� �q�b��q����q7� ���`�گ����� ��*��؟R�� �z� �(����P�ʿ�x� ������ȯB�D� ���r�p��p���� <��������	�B�-� f�Qߊߜ߇��߫��� �����,��>�b�M� ��q��������� ��(��L�7�p�[��� ������������� 6!ZlW�{� �����2�V�z_DEV ���MC:���T4��pGRP 2�����p�bx 	� 
 ,�^��� �/�&///\/C/ �/g/�/�/�/�/�/�/ ?�/4??X?j?��? E?�?�?�?�?�?OO OBO)OfOMO_O�O�O �O�O�O�O�O_q?_ P__t_[_�_�_�_�_ �_�_o�_(ooLo^o Eo�oio�o�o�o�o3_  �o6ZAS �w������ �2�D�+�h�O����� �oy����ߏ�� @�R�9�v�]������� П����۟�*��N� ��C���;�����̯ޯ ů��&�8��\�C� ����y�����ڿ��ӿ �g�4�F�-�j�Qώ� uχ��ϫ������� �B�)�f�x�_ߜ߃� ����)��߭��,�� P�7�t��m����� �������(��L�^� E�����w���o�����  ��6ZlS �w�����p�D��d Ԗ�	2{f������O%��/�����4!�4%D/R' </r/`/�/�/�/�)/ �/0)�/??>?,?N? P?b?�?�/�?�/�?�? �?OO:O(OJO�?�? �O�?pO�O�O�O�O_  _6_xO]_�O&_�_"_ �_�_�_�_�_oP_5o t_�_hoVo�ozo�o�o �o�o(oLo�o@. dR�v�� � $���<�*�`�N� �������t���p�ޏ ��8�&�\����� L�����Ɵȟڟ��� 4�v�[���$���|��� ��¯į֯�N�3�r� ��f�T���x������� �:��J��>�,�b� Pφ�tϪ����Ϛ� ߖ��:�(�^�L߂� �ϩ���r����� ��� �6�$�Z�߁���J� ������������2� t�Y���"���z����� ������:�1��
 ��R�v��� �6�*:<N �r����/ �&//6/8/J/�/� �/�p/�/�/�/�/"? ?2?�/�/?�/X?�? �?�?�?�?�?O`?EO �?OxO
O�O�O�O�O �O�O8O_\O�OP_>_ t_b_�_�_�_�__�_ 4_�_(ooLo:opo^o �o�o�_�oo�o �o $H6l�o�� \~X��� �� D��k��4������� ������^�C��� �v�d����������� ��6��Z��N�<�r� `���������"��2� ̯&��J�8�n�\��� ԯ�������~���"� �F�4�jϬ���пZ� �ϲ���������B� ��iߨ�2ߜߊ��߮� �������\�A��
� t�b�������"� ��������:�p�^� �������������  "$6lZ��� �������  2h���X� ���
/�/p� g/�@/�/�/�/�/�/ �/?H/-?l/�/`?�/ p?�?�?�?�?�? ?O D?�?8O&O\OJOlO�O �O�O�?�OO�O_�O 4_"_X_F_h_�_�O�_ �O~_�_�_o�_0oo To�_{o�oDofo@o�o �o�o�o,noS�o �t����� �F+�j�^�L��� p�������܏��B� ̏6�$�Z�H�~�l��� �
�۟������2�  �V�D�z�������j� ԯf��
���.��R� ��y���B�����п�� ����*�l�Qϐ�� ��rϨϖ��Ϻ���� D�)�h���\�J߀�n� �ߒ���
������� ��"�X�F�|�j���� ��������
��� T�B�x������h��� ������P�� w��@����� �X~O�(� p�����0/ T�H/�X/~/l/�/ �/�//�/,/�/ ?? D?2?T?z?h?�?�/�? ?�?�?�?O
O@O.O POvO�?�O�?fO�O�O �O�O__<_~Oc_u_ ,_N_(_�_�_�_�_�_ oV_;oz_ono\o~o �o�o�o�o�o.oRo �oF4jXz|� ��*���B� 0�f�T�v���Ï� �������>�,�b� ����ȏR���N�̟� ����:�|�a���*� ��������ȯ�ܯ� T�9�x��l�Z���~� ����Ŀ�,��P�ڿ D�2�h�Vό�zϰ�� ���Ϡ��Ϝ�
�@�.� d�R߈��ϯ���x��� �������<�*�`�� ����P��������� ���8�z�_���(��� ������������@�f� 7v�jX�|� ���<�0� @fT�x��� �/�,//</b/ P/�/��/�v/�/�/ ?�/(??8?^?�/�? �/N?�?�?�?�? O�? $Of?KO]OO6OO~O �O�O�O�O�O>O#_bO �OV_D_f_h_z_�_�_ �__�_:_�_.ooRo @obodovo�o�_�oo �o�o*N<^ �o�o��o���� �&��J��q��:� ��6���ڏȏ���"� d�I����|�j����� ��֟ğ��<�!�`�� T�B�x�f�������ү ���8�¯,��P�>� t�b���گ��ѿ���� ���(��L�:�pϲ� ��ֿ`��ϸ������� $��Hߊ�o߮�8ߢ� ���ߴ������� �b� G���z�h����� ����(�N��^���R� @�v�d������� ��� $�����(N<r `��������� $J8n�� �^����/�  /F/�m/�6/�/�/ �/�/�/�/?N/3?E? �/?�/f?�?�?�?�?��?&?OJ?L1�$S�ERV_MAILW  T5J@�0H�OUTPUT?H�0HRV �2��6  M@ �(�1O�O4DTOP�10 2�I d P?�O�O__ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9K] o�������5ιEYPE`LNEFZ�N_CFG ��5MCL4oB�?GRP 2�%��� ,B   A�e�L1D;� B�f��  B4L3�RB21�FHELL���5��@�O<�ΏK%RSRݏޏ��)��M� 8�q�\�������˟����ڟ���7�I�[��  �+�[���X��i��� L0��PŢơL8q�2L0d��������HK 1��� ˯@�J�D� n���������߿ڿ� ��'�"�4�F�o�j�|���ϊ�OMM �����Ϗ�FTOV_�ENB?D�A��O�W_REG_UI���2BIMIOFW�DL�����h�3�WAIT����oE^��Z@��DX�TIMn�����VA>@|i�3�_UNIT������LC�TRY���4@MON�_ALIAS ?5e���@heOM� _�q��J;������ ���� �2�D�V�� z���������m����� 
.��Rdv� 3������ *<N`��� ��w�//&/8/ �\/n/�/�/=/�/�/ �/�/�/�/"?4?F?X? j??�?�?�?�?�?�? �?OO0O�?AOfOxO �O�OGO�O�O�O�O_ �O,_>_P_b_t__�_ �_�_�_�_�_oo(o :o�_^opo�o�o�oQo �o�o�o �o6H Zl~)���� ��� �2�D��h� z�������[�ԏ��� 
��Ǐ@�R�d�v��� 3�����П⟍��� *�<�N���r������� ��e�ޯ���&�ѯ J�\�n���+�����ȿ ڿ쿗��"�4�F�X� �|ώϠϲ���o��� ����0���T�f�x� ��5߮��������ߡ���,�>�P�b���$�SMON_DEF�PROG &������� &*SYST�EM*i�����<{�RECA�LL ?}�� �( �}3xco�py fr:\*�.* virt:�\tmpback���=>192.1�68.56.1:?17836 � �X2�D��}4��a������������ }�8��s:orde�rfil.dat�v�����/AS}/��mdb:s�� ���`���z�� �.@Re���� �������~�*/ </N/as/��/�/ �/�r�&?8?J? ]o ?��?�?�?� �v//"O4OFOY/k/ O�/�O�O�O�/�/|? ?�O0_B_�Og?�O
_ _�_�_�_�?�?�O�O ,o>oPocO�_�Oo�o �o�o�Ot_�__(: L__�o�_��� �_�_xoo$�6�H�[o mo��o����Ə�o�o ~ �2�D�Wi�� ����U����� ��.�@�R�e� ���� ����Я�v����*� <�N�a��������� ̿ߟ�z��&�8�J� ]�o�
ϓ��϶���ۯ ���"�4�F�Y�k� �Ϗ��߲���׿��� �ߟ�0�B���g��� ��������x߅�� ,�>�P�c�����ߪ� ��������|��(: L_�s����� ������$6H[� m����������� t� /2/D/Wi/��/�/�/U.�$S�NPX_ASG �2�����!��  0��%��/?  ?���&PARAM ���%�! ��		;P����o4�� OFT�_KB_CFG � ��%�#OPI�N_SIM  
�+j2�?�?�?�3�� RVNORDY?_DO  t5�5�BQSTP_D�SB�>j2HO�+S�R ��) �� &n:�O��&T�OP_ON_ER�RO�FPTN ��%�@�C��BRING_PR�M�O#BVCNT_�GP 2��%l1 0x 	DO?_�-_�f_Q_�_�'VDPROP 1�C9m0{Q �1m_�_�_�_�_o4o 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu����� ����)�;�M�_� ����������ˏݏ� ��%�L�I�[�m�� ������ǟٟ��� !�3�E�W�i�{����� ��دկ�����/� A�S�e�w��������� ѿ�����+�=�d� a�sυϗϩϻ����� ���*�'�9�K�]�o� �ߓߥ߷��������� �#�5�G�Y�k�}�� ������������� 1�C�U�|�y������� ��������	B?�Qcu���RPRG_COUNT�6s��B�	ENB�O��M��4�_UP�D 1�nKT  
��ASe� �������/ /+/=/f/a/s/�/�/ �/�/�/�/�/??>? 9?K?]?�?�?�?�?�? �?�?�?OO#O5O^O YOkO}O�O�O�O�O�O �O�O_6_1_C_U_~_ y_�_�_�_�_�_�_o 	oo-oVoQocouo�o �o�o�o�o�o�o. );Mvq��� ������%�N� I�[�m���������ޏ�ُ돷_INFOg 1�/ �� �R�=�v�a���������YSDEBU)G� 0���d��SP_PASS��B?�LOG ��/9  ������  ����UD1:�\�ϟ �_MPC $�/����/[�Я� /��SAV ��'����G�_����f�SVԛTEM�_TIME 1��'�: 0  ����W�f�ўTSKMEM  /��G�  ��%ps���Ͽ��� @���� �������U��A������J�*\�n�(�����ϐ�ϸ���^��� W����p�+�=� O�a�s߅ߗߩ߻���������u�9�K� ]�o��������� �����#�5�G�Y�k��}���T1SVGgUNS*�'����ASK_OPTION� /���_DI�����BC2_GRP �2�/�Q�%��@��  C�:��BCCFG ��� ����` ��������! E0iT�x� ����/�/// ?/e/P/�/t/�/�/�/�/�/?���,!?�/ T?f?�/C?�?�?�?�? �?׮O���0O2O O VODOzOhO�O�O�O�O �O�O�O_
_@_._d_ R_t_�_�_�_�_�_�_ o�_oo*o`oFh10 to�o�o�o�oFo�o�o �o"FXj8� |������� 0��T�B�x�f����� ��ҏ�������>� ,�N�P�b�������ro ԟ���(���L�:� \���p�����ʯ��� ܯ� �6�$�F�H�Z� ��~�����ؿƿ��� �2� �V�D�z�hϞ� �Ϯϰ��������ҟ 4�F�d�v߈�߬ߚ� ��������*���N� <�r�`������ ������8�&�\�J� l��������������� ��"XF|2� �����f� B0fx�X� �����/// P/>/t/b/�/�/�/�/ �/�/�/??:?(?^? L?n?p?�?�?�?�?� �?O$O6OHO�?lOZO |O�O�O�O�O�O�O_ �O2_ _V_D_f_h_z_ �_�_�_�_�_�_o
o ,oRo@ovodo�o�o�o �o�o�o�o<�? Tf���&�� ���&�8�J��n� \���������Əȏڏ ���4�"�X�F�|�j� ������֟ğ���� �.�0�B�x�f���R ��Ư������,���<�b�P���p���A���*SYSTEM�*��V9.005�5 ��1/31/�2017 A �v  ��K�T�BCSG_GRP�_T   \ �$ENABLE��$APPRC�_SCL   
$OPEN��CLOSE�S_�MINF2'�AC�C��PARAM�� ���MC_MAX_TRQ�{$d�_MGNk��C�AVw�STA�Lw�BRKw�NO�LDw�SHORT?MO_LIM�ʧ�rh�J����PL1��T6���3��4��5��6��7��8k�s��~�� $DъE�E��T��b�P�ATH^�w�m�w�_RATIOk�s�T�� 2 	$CNT�A�����m�{INX�_UCA����CAT_UM���YC_ID 3	����_E�����6������PAYL�OA��J2L_U�PR_ANG6�L�WA�?�3�O�x�R_F2LSHRTv�LOD���}��Ӌ���?ACRL_S�ؽ���+�k�HVA��$Hx���FLEX�� �J2�� P�B_F���$��_FTM���&��$RESECRV�>�;������� :$���LEN.�z�;�DE|���;�Yғؔ���SLOW_AXI^��$F1��I���2��1������MO�VE_TIM��_?INERTI��
��	$DTORQCUEX�3��#I��ACEMN��%E�%Ep	V��d�A8�R�TCV��@Rt����
��T@�RJ���	�M��,��J_�MOD����� �dRy�2��P�pE���\�X���AW�gQJKh@��K��VK�;VK�JJ0����JJ�JJ�AA6��AA�AA%�3AA �t�N1�N �d�#��E_NUv�� �CFG�� � $GR�OUPc�SK��B�_CON�C��B�_REQUIRE����BU��UPD�ATT�EL�}  �%� $kTJ��� JE��gCTR��
TN �F�&�'HAND_kVB��OP�7 $oF2x�3��m�COMP_SW������R��� $$Ma�e�R �Î8���<� �5�¼6�A_.�h�D�<q�A*��A��A��A���0���D��D��D��Pf��GR�ǂAST��h�A�ɂAN��DY�� �x��4�5A���s�� s��2�B��R����P����� �)��2�;�s2J� �0i�\� 7�U6���QASYM��
��TС��мݎ���_SH�"�������TU8 ����%�7�J>����P�pcfio�_VI�83�h6þ`V_UCNI���d�{�JU �bU�b���d���d v ����������su���� �r2�HR_T��	N2�q���DI����O�tr2�pN�#
  �2I�QAz����q �S�s �� � �p  �� f1MEeМ��pr�QT�pPT@&`r a�>���~$�5`C�^�R�T4`!� $DUMMY}1�$PS_ �RF��$��n��FLA� YP_���F�$GLB_T�0�u΅>���t0; 1�q X��'��STf� SBR�v�M21_VT�$SV_ERa�O�(`�,�CL��A�p O�r�pGL�`E�W� 4 $�H�$Y�2Z�2Ww��x�b3A����Y�U]� oN���)`$GI0{}$]� �q8Z���� Lh����'b}$F'bE��NWEAR_ N��F��\ TANC�Ҥ���JOG���� �e�$JOINT�& f�Y�MSET.�  ��E�« S�✔�!�׼  Ue?��� LOCK_FOx��m1�pBGLV3�GL��TEST_sXM�j�EMP=��Ϣ悖�$UC�\���2� �������i0�����C�E| Ó� $KA�R�M�sTPDRqA`�3�*�VEC~��D�.�IU���!CH=E��TOOL��i��V��REK�IS3�;���6���ACHP���v�O��F����29���I�� � @$RAIL_�BOXE�� R�OBOƤ?��HOWWAR��屖���ROLM���q!���¡!Ӱ��J�O_=F� ! �!Y����K�6�=0RN�OBo�6���?�C��s�Z�OUR������Q�"�!��$PIPǦN]�Ӳ�� ���V�@�CORDEAD����u��p� O�p  D ̀OBA�#�������p̀��'`�!SYS���ADR�!�p>�TC}H�0  ,oSEN�r#�A��_���d�z!�ћrVWV�A� � �9�]��uPREV_�RTA$EDI}T��VSHWR�!��&��]q��`D�(�.Q��6Q$H�EAD8amp��Ha��KEq�|�CPS�PD�JMP�Ld�ut0Ra �t��T�\�IРS�"C20�NEr��!�'TIC�K���QM�QjR:�H=N�� @�W�~%�_GP��ʶ$�gSTY^ү�LO��q3:��� t 5
��Gj�%$�Ѳ�u=��S�!$�a Jp-����p��P�P��SQU-������aTGERCB�gQt0S�$ ����']�'-`�>pOC�6�bP�IZ��������P�R������S��PU��a��_DO�c�XuSN�K�vAXI��/���UR� p�" 찕�"�]1� _`�4ҋET5P��ЦU���F�W��A�A�Q���ĳ��!r2S=RE4lu��9 ��:��6�	�2��7 ��9��9�G�G �'F"TIF�R&��4CE o2o�DoVdU�SSCЀ o h� DS���4���SP�p"%AT�@�2���c⅂A_DDRESs�B���SHIF�#�_2+CH� �I�t!��TU�I�1 }6�CUSTOV*�V��I�r UҸ��6!��P
Ϫ
�V8������! \����A����,��J�2CSC���Y�*��2�1�T�XSCREE��"z�p�TINAO�x��T4��  *j�sQ_6"vP# TI� /���4�.���63�8�4��RRO�@�`3�
��1F�UE?�G$ ��PMѧ�SP��4�RSM����UN�EX_�vA�pS_ ��+F�SA.IIG�S6�C��B�4 2#O0UErT%�r?�nF���GMT3pL�a��O@�kPBBL�_��Wo���& �����BO���BLE�f"�C밚"�DRIG�H�CBRDA�\!C�KGRo�UTEX�$ UQWIDTH@����Ʊ��Jq�0�I>�EY6 ��' Adh�0�����Ӱ��BACK�ᡂ�UE��!�FO���WLA-B�?(!�I����$UR��P�@_P�'�H�1 ( 8�wq�_��t"�R(�R�q�����������QO�m!��)��L�PU��@7cR���LUM87cV ERV��U�R_PP�fT*�j CGE�R�a `�)��LP�e_E\���)��g��h!�h���i5*�k6�k7�k8�bZ�@6����4�������SJ�)^QUSR�]�+ <��'�U����#��FO� ��P�RIrm��%q�pT�RIPϱm�U)N�p�t,����p�����/��3 -� q-�RSp��G  �aT/��u!�rOSF���vR9 �2�so���.`f�x����� �s	U�a��/$�6�DC�b����sOFFŠ��0���L�O�� 1�.9�����/9�GU.�P���׃��sQ�SUB��H��@SR	T��1���;���sOR��'�RAU� r(�T=�Z��VC� >Ҕ2� ɲ���$���y�8񹳬`C���{�DRIV���@_V�����Ѐ�D~4tMY_UBY3t �����$��19�l0��q	����P_S������BM�A$nb�DEY_�EX�@��3����_MU.�X�An� @US2�8��p�[�k0w�xp� �2x�G>gPACINr�!�RG�𦥽�����A���SCp�RE�Rj!o��`���S�3 ^Y�TARGÐP72H��a�R�S�4nP�0`TQ�	o���RmEz�SW��_A���� o���OIq\!A(n v��E$pU�෱�� �0a�HK��5����W�s��0��sEA��ɷWOR�Pxv��0�MRCV�AW6 ��`O��M�P�C83	����REF�G(����e�s` cM�Xp�^��^�-�8��Ƶ�_RCʻ���0S!pf�ϓ��L8~@`��D7 ���gP�TU0 epԕw�OU�����惓 2��2 $U00��Fr�45#�^�K �SULg 5c`CO�0 `6`�]��� �0���Ѫ�a��@q��i�L���$���a���@q�s�?�8|� +5#k� 5#C7ACH��LOR�&��<�a�A�KQC ��C_oLIMIg#FRj�qTl���$HO�Pz�*�COMM��BO�@��ب �a�F�VP��/ ��_�����Z����k���WAv{�MP�FAIk�5G��;�AD?�p��IMRE�_���G�P@V�� k�ASY�NBUFk�VRTaD������&SOLo SD_|���WA�P�'ETUO�X�Q�����ECCU�VEM�٠%�k�VIRC�?����B��_DE�LA����p�p�AuG��Rc�XYZM@�5Cc�W3�qsQ T ��P�[Qs��D9�"�Q�LASAP�
�� G$l� :�rX�Sa�7��N�m�VLEXEE�;�3W�ka5!�y�FLPIW���F�I����F���P�q9#�<_p�
���8t@s���@ORDB|q���##�� =_0�Z`T�r�B�O|JP6b�VSFE �3>  a0s���c��UR� �SM�u�?�rV�R J� f��"�5@�r��qgLIN��@�WN�XS屎 A��2��uK&SHd`HOLk��P�XVR�tB|��@T_OVRk� �ZABC�C ��"q-1
�Zހ�t}D�rDBGLV���Lϒ�R]�ZMP�CF�E�0�t�2ޑLN~ ��
81d��F Ђ`��ɰ4CMCM��C>��CART_Y1���P_2` $	Jw3q4D��}2�2�70`�5`��UX|5�UXEu��6|�5��4�5�1�1�9�1�6
y� �%G +T�$��CBYV D�p H�RRM�{q��CHET����PU'�Q�!P�I �� ��A� PEA�Kf���K_SHIX�B��'RV F^`G½B� C�@r2g1|� ����A20��I S��}DXTRACE�P�V�"ASPHER'aJ ,e�THjO�|I��$TBCS�G� 2 ��}��Q���}��   
 ` �_�_�_�_�_�_�_��_.ooRodkwR~S~�\d ��a}?�Q	 HCBdo~�iC  B �R0�o�h�o�kB��o�p��o�jdf  AXp?�w{qW� {������@�@� :nT�g�z�E�W� �������
����3�	V3.0�0�R	md45N�	*U�M����1�� ��m����  ��֟�wQJ2{c�]6���� � �U�Q ,����E�şp�G�p�����	_� ȯ���ׯ���4�� D�j�U���y�����ֿ �������0��T�?� x�cϜχϬ��Ͻ���@����>�P�X�7� j�|�&ߜ��߬����� 	���-��Q�c�u�� B���������� �U%�7��Q��=�c�Q� ��u������������� ��)M;q_� ������ 7%GI[�� �������// �M/;/]/�/q/�/�/ �/�/�/??%?�/I? 7?m?[?}?�?�?�?�? �?�?�?!OOEO3OiO WOyO�O�O�O�O�O�O _�O__/_e_S_�_ w_�_�_�_�_�_o�_ +ooOo=oso�o//�o �o5/ko�o�o9 'Io]���u �����5�G�Y� k�%���}�������� ׏���1��U�C�e� ��y�����ӟ����� �	��Q�?�u�c��� ������ͯ����o �oA�S���+�q����� ��ݿ˿��%�7�I� [���mϏϑϣ��� �������3�!�W�E� {�iߋߍߟ������� ����A�/�Q�w�e� ������������� �=�+�a�O���s��� ��e���������' K9[]o��� ����#G5 k}��[��� ��//C/1/g/U/ w/y/�/�/�/�/�/	? �/-??=?c?Q?�?u? �?�?�?�?�?�?�?)O OMO_O��wO�O3OaO �O�O�O�O__7_%_ G_m__�_O_�_�_�_ �_�_o!o3oEo�_io Wo�o{o�o�o�o�o�o �o/SAce w������� �)�O�=�s�a����� ����ˏ�O	��-� ׏]�K���o������� ۟ɟ���#�5��Y� G�}�k�����ůׯ�� ����1��U�C�y� g�������ӿ����� �	�?�-�O�Q�cϙ� �Ͻϫ��������� ;�)�_�M߃ߕ�?��� ��i������%��I� 7�m�[�}������������!��E�/� s e�i� i��}�i��$TBJO�P_GRP 2�1�� / ?�i�	�������9� ?� ����+ ��������i�� @e��	 ��CB  ��C�����5GU	i�C� 2BH  A��/��D�,��bB* q��$�7C��  ���c�d�L�i�A �EG+ ��a	���D/�D<Ky/�//#/�/�/��	??�/�/ T?f?%?o?a	�?�?�? �?�?�?�?O)OO!O OO�O[OO�O�O�O�O(�O_g�i�1Q�E	V3.00���md45��*�[P��d�i_tW �G/� G7� �G?h GG8 �GO Gd� �Gz  G�� �G�| G�: �G�� G�� �G�t G�2 �G�� Gݮ �G�l G�* G�� HS�R�F� F@ �F+� FK  �Fj` F� �F�Q � GX� �R�Q^� Gv� G�ĨS�4� G�� G��� G�\ G�� =L��=#�%
]Ae�Js�Yo�kbi�oo�o��E_STPAR�P]����HR�`ABL�E 1	��C`i��h�g ��di�g��hn i�h�p�g	��h
�h�h�ei���h�h�hDa�cRDI�o���o!3EWu�tO��{� ���+��bS��� �z����"�4�F� X�j�|�������ğ֟ �����0�B���Ā ȏ���g��l�~����� N`r���x�bi��NUM  1�U��	 q� C`�D`�b_CFG �
R���@��IM?EBF_TT�a��8���`��VERBc��z����R 1�kO 8f_i�d�2� 4���  �� �%�7�I�[�m�ϑ� �ϵ����������!� 3�|�W�i߲ߍߟߵ�������A�����cMD3�E��� k�}��V_I����GINT�����T1�#�5� B��O�a���G_TC������$�P����9�RQ��Դ�_L���@˵�`M�I_CHAN�� �˵ nDBGLV�L��˵�aq ET�HERAD ?*�e� ��`������hq ROUT6��!P�!#A~SNMASK�|˳�255.�GS}��GS�`OOLOFS_DI�P��%�	ORQCTRL ޻7��o-T/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?s</�?�?��?�cPE_DET�AI��PGL_�CONFIG �R�b���/c�ell/$CID?$/grp1�?4O FOXOjO|O2��
�O �O�O�O�O_�O%_7_ I_[_m___�_�_�_ �_�_�_�_�_3oEoWo io{o�oo�o�o�o�o �o�o/ASew �*��������}�O�a�s���@������?я���� ��*�<�N�`���� ������̟ޟm��� &�8�J�\�n������� ��ȯگ�{��"�4� F�X�j���������Ŀ ֿ������0�B�T� f�x�ϜϮ������� �υ��,�>�P�b�t� ��ߪ߼�������� ��(�:�L�^�p��� ��������� ��@��User �View "I}}�1234567890C�U�g�y��������. C����)�2 6���+=Oa����0�3�����@��	h*��4� cu�������5R/)/;/M/_/q/��/��6/�/�/��/??%?�/F?��7 �/?�?�?�?�?�?8?�?��8n?3OEOWOiO�{O�O�?�O�B �lCamera4�*O�O__)_;_M_+�E�Ow_�_�^A���_�_�_�_�_o)  �F���O_oqo�o�o �o�o`_�o�oLo%@7I[m�O��F �	�����%� �oI�[�m�������� Ǐُ돒�wQ��7� I�[�m����8���ǟ ٟ$����!�3�E�W� ���w+k🥯��ɯۯ �����#�5�G���k� }�������ſl��E�) Z��!�3�E�W�i�� �ϟϱ���������� �/�ֿ�wm9��{ߍ� �߱�����|����� h�A�S�e�w���B� �w!I2�������/� A���e�w��������@����������9�� HZl~��I�� ����� 2DV(hz	J	�E0 � ����/�3/E/ W/�{/�/�/�/�/�/ |��@�Ky/.?@?R? d?v?�?//�?�?�?? �?OO*O<ONO�/�E Bk�?�O�O�O�O�O�O �?_*_<_�O`_r_�_ �_�_�_aO��{Q_o o*o<oNo`o_�o�o �o�_�o�o�o& �_�U��or��� ��so���_8� J�\�n�����9�U�� )�ޏ����&�8�� \�n���ˏ����ȟڟ ������U򻕟J�\� n�������K�ȯگ� 7��"�4�F�X�j��  ������� Ͽ����)�;�M�_�   o�w��� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e��w�����������c� � 
�(  �>��( 	 �� ;)_M�q� �����%��� ̹�j| �������/ �Y6/H/Z/�~/�/ �/�/�/�//�/? ? g/D?V?h?z?�?�?�/ �?�?�?-?
OO.O@O ROdO�?�?�O�O�OO �O�O__*_<_�O`_ r_�_�O�_�_�_�_�_ oI_&o8oJo�_no�o �o�o�o�oo!o�o "ioFXj|�� �o���/��0� B�T�f��������� ҏ�����,�s��� b�t���͏����Ο�� ��K�(�:�L���p� ��������ʯ�� � �Y�6�H�Z�l�~��� ׯ�ƿؿ�1�� � 2�D�V�hϯ��Ϟϰ� ��������
��.�u� R�d�v߽Ϛ߬߾���p����;�@ �#�5�G��� ���0frh:\t�pgl\robo�ts\am100�id\arc_m�ate_��_14?50.xml�� ����������0�B�T�E���Y�~����� ���������� 2 D[�Uz���� ���
.@W Qv������ �//*/</SM/r/ �/�/�/�/�/�/�/? ?&?8?O/I?n?�?�? �?�?�?�?�?�?O"O 4OK?EOjO|O�O�O�O �O�O�O�O__0_GO A_f_x_�_�_�_�_�_��_�_oo,o>n`�Ζ� �k�<<w i�?�>k �o>oyo�o�o�o�o�o �o�o5-O}c ���������1�?��$TPGL�_OUTPUT �I�I� a`i�~������� Ə؏���� �2�D� V�h�z�������ԟ@���
��i�a`�6��2345678901A�S�e�w����� ��?�>�ʯܯ� �� $���(�Z�l�~�����:�}��Կ���
�� ��ƿR�d�vψϚϬ� DϺ�������*��� 8�`�r߄ߖߨ�@�R� ������&�8���F� n�����N����� ���"�4�����j�|� ��������\����� 0B��Px�� ��Xj�, >P�^���� �f�//(/:/L/�A�}\a�/�/�/�/�/�/�-@co?#?ij ( 	 &� X?F?|?j?�?�?�?�? �?�?�?OOBO0OfO TO�OxO�O�O�O�O�O _�O,__<_>_P_�_t_�_4��_`xf�_�_ �]�_o*ooNo`o.� �_�o�o=o�o�o�o�o !o%W�oC� �y��3��� �A�S�-�w����q� ��яk������=� ����s���������� ����a�'�9�ӟ%� o�I�[��������� ��ٯ#�5��Y�k�ɯ S�����M�׿�ÿ� �}��U�g�ϋϝ� wω���1�C�	�ߵ� '�Q�+�=߇ߙ��ϝ� ��i߻�����;�M� ��5���o����� ���_���7�I���m� �Y������%����� ��3i{�� ��K�����/�R�$TPOF?F_LIM �P�>�Q��J�N_SVN  ��$`P_MON7 �Ub���2�%JSTRTCHK �U�`/hVTCO�MPATu�dVWVAR ��"(y � �:/Y�J_D�EFPROG �%�%Q/�/f_DISPLAYU��j"INST_M�SK  �, ~�*INUSER�ά$LCK�,�+QU?ICKMEN"?�$oSCREA0�U~ "tpsc�$��!\0a9`r0_v9S�T�`RACE_�CFG ��"$Y	C$
?�~�8HNL 2y*�P�1)+ O"O'O9O�KO]OoO�O�O�J�5I�TEM 2K� �%$1234?567890�O�E  =<�O_*_2S�  !8_@[L  �O�_C#�O�_
_�_�_ @_�_d_v_?o�_Zo�_ jo�oooo*oDoNo �oroDV�oz�o �o|&��
�n ����:������ ��"�ʏF�X�!�|�<� ��`�r�֏����L�՟ 0��T� �&�8���D� ��ҟ�^����گ� P��t������4�ί �������(�:��^� ς�B�Tϸ�j�ܿ� �����6���ߎ�~� �Ϣϼ���@��ϖ߼� ��2���V�h�z��ߞ� J�p���ߎ�
��.� �� �d�$�6���B��� �����������N�  r���M��h��x ���8J\� �,Rd���� ��F//|$/ ��{/��/��/�/@0/�/T/f//?�4S�2��?4:�  ��B4: �1�?�)
� �?�?�?�?c:�UD1:\�<���F1R_GRP 1��K� 	 @� :OLK6OlOZO�O~O�O�N��@�O�J��A�?_�O7_"U?�  R_d[N_�_r_�_ �_�_�_�_�_�_&oo Jo8ono\o�o�o�o�o�	5�o�oD3SC�B 2P;  =_:L^p������:<UTORIAL P;�?��?7V_CONFIG  P=�1�?�?�t�$�OUTPUT� !P9e�����ď֏����� 0�B�T�f�x�����b� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���(�:�L�^�p� �ϔϦϷ������� � �$�6�H�Z�l�~ߐ� �߳���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r�������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/N�`����/??&? 8?J?\?n?�?�?�?�? �?��?�?O"O4OFO XOjO|O�O�O�O�O�? �O�O__0_B_T_f_ x_�_�_�_�_�_�O�_ oo,o>oPoboto�o �o�o�o�o�_�o (:L^p��� ���o� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶�����Ͻ(��� �������6��/Z�l� ~ߐߢߴ��������� � �2��V�h�z�� �����������
�� .�@�Q�d�v������� ��������*< M�`r����� ��&8I\ n������� �/"/4/F/Wj/|/ �/�/�/�/�/�/�/? ?0?B?S/f?x?�?�? �?�?�?�?�?OO,O >OO?bOtO�O�O�O�O �O�O�O__(_:_L_ ]Op_�_�_�_�_�_�_ �_ oo$o6oHoY_lo ~o�o�o�o�o�o�o�o� 2DS{�$T�X_SCREEN� 1"����}�S�������Bք 1�C�U�g�y����� ��ӏ���	����?� ��c�u���������4� �X���)�;�M�_� ֟蟕�����˯ݯ� f����7�I�[�m�� �����,�ٿ���� !�3Ϫ���i�{ύϟ� ����:���^���/��A�S�e��ω��$U�ALRM_MSG� ?sy��p  ��Vj��������"�� F�9�K�i�o�����������SEV  ������EC�FG $su�}q  Ve@� � AJ�   B�Vd
 ��]csu}� ���������������1?&�GRP �2%0� 0Vf	� g����I_B�BL_NOTE �&0�T�G�l]bxp_a<�~�DEFPRO��<Z�� (%�� _`�*N9r] �������/��FKEYDAT�A 1'sys ps ?�Vf =�x/�/� g/�/�/�%,(/�/Vd�/??C? *?g?y?`?�?�?�?�? �?�?�?O-OOQO8O uO�OnO�O�O�O�O�O0_�O)_X.��9_`_ r_�_�_�_�_]bN_�_ �_oo+o=o�_aoso �o�o�o�oJo�o�o '9K�oo�� ���X���#� 5�G��k�}������� ŏ׏f�����1�C� U��y���������ӟ b���	��-�?�Q�c� 򟇯������ϯ�p� ��)�;�M�_�� ������˿ݿ�~�� %�7�I�[�m�D_�ϣ� ����������!�3� E�W�i�{�
ߟ߱��� �����߈��/�A�S� e�w��������� �����+�=�O�a�s� ������������� ��'9K]o�� "������ 5GYk}�� ����//�C/ U/g/y/�/�/,/�/�/ �/�/	??�/??Q?c?�u?�?�?�?���;}�������?@�?�=�? O2OF,_ cO_�OnO�O�O�O�O �O__�O;_"___q_ X_�_|_�_�_�_�_�_ o�_7oIo0omoTo�o �o���o�o�o�o! 0?EWi{��� @�����/�� S�e�w�������<�я �����+�=�̏a� s���������J�ߟ� ��'�9�ȟ]�o��� ������ɯX����� #�5�G�֯k�}����� ��ſT������1� C�U��yϋϝϯ��� ��b���	��-�?�Q� ��u߇ߙ߽߫����� �o��)�;�M�_�f� �����������~� �%�7�I�[�m���� ����������z�! 3EWi{
�� �����/A Sew���� ��/�+/=/O/a/ s/�//�/�/�/�/�/ ?�/'?9?K?]?o?�? �?"?�?�?�?�?�?O �?5OGOYOkO}O�OO �O�O�O�O�O__���![������J_\_n]F_�_�_|V,�o�_�o�_�_o -ooQo8ouo�ono�o �o�o�o�o�o); "_F�j��� ������7�I�[� m�����O��Ǐُ� ���!���E�W�i�{� ����.�ß՟���� ���A�S�e�w����� ��<�ѯ�����+� ��O�a�s�������8� Ϳ߿���'�9�ȿ ]�oρϓϥϷ�F��� �����#�5���Y�k� }ߏߡ߳���T����� ��1�C���g�y�� �����P�����	�� -�?�Q�(�u������� ��������); M_������� �l%7I[ ������� z/!/3/E/W/i/� �/�/�/�/�/�/v/? ?/?A?S?e?w??�? �?�?�?�?�?�?O+O =OOOaOsOO�O�O�O �O�O�O_�O'_9_K_ ]_o_�__�_�_�_�_ �_�_�_#o5oGoYokoh}o�of��k�f�����o�o�m�o �f,�C� gN������ ����?�Q�8�u� \�������Ϗ���ڏ �)��M�4�q���b� ����˟ݟ��o%� 7�I�[�m���� ��� ǯٯ������3�E� W�i�{������ÿտ ����Ϭ�A�S�e� wωϛ�*Ͽ������� �ߨ�=�O�a�s߅� �ߩ�8��������� '��K�]�o���� 4����������#�5� ��Y�k�}�������B� ������1��U gy������� �	-?Fcu �����^�/ /)/;/M/�q/�/�/ �/�/�/Z/�/??%? 7?I?[?�/?�?�?�? �?�?h?�?O!O3OEO WO�?{O�O�O�O�O�O �OvO__/_A_S_e_ �O�_�_�_�_�_�_r_ oo+o=oOoaosoo �o�o�o�o�o�o�o '9K]o�o��@������ ���� ����*�<�N�&�p���\�, n���f�׏������ 1��U�g�N���r��� �����̟	���?� &�c�J����������� ����)�;�M�_� q��������˿ݿ� ϐ�%�7�I�[�m�� ϣϵ��������ό� !�3�E�W�i�{ߍ�� ������������/� A�S�e�w����� ����������=�O� a�s�����&������� ����9K]o ���4���� #�GYk}� �0����// 1/�U/g/y/�/�/�/ ��/�/�/	??-??? �/c?u?�?�?�?�?L? �?�?OO)O;O�?_O qO�O�O�O�O�OZO�O __%_7_I_�Om__ �_�_�_�_V_�_�_o !o3oEoWo�_{o�o�o �o�o�odo�o/ AS�ow���� ��r��+�=�O� a����������͏ߏ n���'�9�K�]�o��F q��F ��������������̖,ޯ#�֯G�.� k�}�d�����ůׯ�� ����1��U�<�y� ��r�����ӿ����	� �-��Q�c�B/�ϙ� �Ͻ���������)� ;�M�_�q� ߕߧ߹� ������~��%�7�I� [�m��ߑ������� �����!�3�E�W�i� {�
������������� ��/ASew� ������ +=Oas�� ����//�9/ K/]/o/�/�/"/�/�/ �/�/�/?�/5?G?Y? k?}?�?�?x��?�?�? �?OO&?COUOgOyO �O�O�O>O�O�O�O	_ _-_�OQ_c_u_�_�_ �_:_�_�_�_oo)o ;o�__oqo�o�o�o�o Ho�o�o%7�o [m����V ���!�3�E��i� {�������ÏR���� ��/�A�S��w��� ������џ`����� +�=�O�ޟs�������л�ͯ߯�0��>�0���
�� .��P�b�<�,Nϓ� FϷ���ۿ�Կ��� 5�G�.�k�RϏϡψ� �Ϭ���������C� *�g�y�`ߝ߄����� �?��	��-�?�Q�`� u���������p� ��)�;�M�_���� ����������l� %7I[m���� ����z!3 EWi����� ����///A/S/ e/w//�/�/�/�/�/ �/�/?+?=?O?a?s? �??�?�?�?�?�?O �?'O9OKO]OoO�OO �O�O�O�O�O�O_�� 5_G_Y_k_}_�_�O�_ �_�_�_�_oo�_Co Uogoyo�o�o,o�o�o �o�o	�o?Qc u���:��� ��)��M�_�q��� ����6�ˏݏ��� %�7�Ə[�m������ ��D�ٟ����!�3� W�i�{�������ï R������/�A�Я e�w���������N�㿀����+�=�O�&P�Q��&P���zόϞ�v����Ϭ�,��߶�'��K�]� D߁�hߥ߷ߞ����� �����5��Y�k�R� ��v���������� ��1�C�"_g�y����� ����п����	- ?Q��u���� �^�);M �q������ l//%/7/I/[/� /�/�/�/�/�/h/�/ ?!?3?E?W?i?�/�? �?�?�?�?�?v?OO /OAOSOeO�?�O�O�O �O�O�O�O�O_+_=_ O_a_s__�_�_�_�_ �_�_�_o'o9oKo]o oo�oX��o�o�o�o�o �oo#5GYk} ������� �1�C�U�g�y���� ����ӏ���	���� ?�Q�c�u�����(��� ϟ������;�M� _�q�������6�˯ݯ ���%���I�[�m� �����2�ǿٿ��� �!�3�¿W�i�{ύ� �ϱ�@��������� /߾�S�e�w߉ߛ߭ߴ�ߖ`����`����������0�B��,.�s�&��� ~����������'� �K�2�o���h����� ����������#
G Y@}d���o� ��1@�Ug y����P�� 	//-/?/�c/u/�/ �/�/�/L/�/�/?? )?;?M?�/q?�?�?�? �?�?Z?�?OO%O7O IO�?mOO�O�O�O�O �OhO�O_!_3_E_W_ �O{_�_�_�_�_�_d_ �_oo/oAoSoeo�_ �o�o�o�o�o�oro +=Oa�o�� �������'� 9�K�]�o�v������ ɏۏ�����#�5�G� Y�k�}������şן ������1�C�U�g� y��������ӯ��� 	���-�?�Q�c�u��� �����Ͽ���� ��;�M�_�qσϕ�$� ���������ߢ�7� I�[�m�ߑߣ�2��� �������!��E�W� i�{���.������������/��$UI�_INUSER � ���P���  �0�4�_MENHI�ST 1(P��  ( �]���(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1o�������� ����936��dv��) ������ ASew��*� ���//�=/O/ a/s/�/�/�/8/�/�/ �/??'?�/K?]?o?�?�?�?�<�D1��D? �?�?OO)O;O>?_O qO�O�O�O�OHO�O�O __%_7_�O�Om__ �_�_�_�_V_�_�_o !o3oEo�_io{o�o�o �o�oRodo�o/ AS�ow���� ��?�?��+�=�O� a�d��������͏ߏ n���'�9�K�]�o� ��������ɟ۟�|� �#�5�G�Y�k����� ����ůׯ������ 1�C�U�g�y������ ��ӿ�����-�?� Q�c�uχϊ��Ͻ��� ����ߔ�)�;�M�_� q߃ߕ�$߹������� ���7�I�[�m�� �� ����������� !���E�W�i�{����� .���������� �Sew����� ���+�� as����J� �//'/9/�]/o/ �/�/�/�/F/X/�/�/ ?#?5?G?�/k?}?�? �?�?�?T?�?�?OO�1OCO.��$UI�_PANEDAT�A 1*����yA  	�}UO�O�O�O�O�O�O )�O_8�O G_Y_k_}_�_�__�_ �_�_�_�_ooCo*o goyo`o�o�o�o�o�o\�o1	� @r /_4FXj|��o �%_�����0� B��f�M���q����� ���ˏ���>�%� b�t�[���|��{C �۟����#�5��� Y��}�������ůׯ >������1��U�g� N���r�����ӿ�̿ 	��-�?ϲ�ğuχ� �ϫϽ���"���f�� )�;�M�_�q߃��ϧ� ���߲������%�� I�[�B��f���� ��L�^��!�3�E�W� i������������� ����A(ew ^������� +O6s���� ������//h 9/��]/o/�/�/�/�/ /�/�/�/?�/5?G? .?k?R?�?v?�?�?�? �?�?OO��UOgO yO�O�O�OO�OF/�O 	__-_?_Q_c_�O�_ n_�_�_�_�_�_o�_ )o;o"o_oFo�o�o|o �o,O>O�o%7 I�om�O��� ���d!��E�W� >�{�b�������Տ�� ����/��S��o�o}�d�������ӟ���)����u�H�Z� l�~�����	�Ư��� ѯ� ��D�+�h�z� a�����¿Կ�����x��c�k�$UI_P�OSTYPE  ��e� �	 �[�*�QU�ICKMEN  �9�H�^�,�RE�STORE 1+��e  '�뿑r�����ϑrm �)�;�M�_� q�ߕߧ߹����߀� ��%�7�I���V�h� z��ߵ���������� !�3�E�W�i�{���� ������������ ��Sew��>� ����+=O as(��� �//'/9/�]/o/ �/�/�/H/�/�/�/�/ ?�?0?B?�/}?�? �?�?�?h?�?�?OO 1OCO�?gOyO�O�O�O�i�SCREy�?�~�u1sc���u2�D3�D4��D5�D6�D7�D8��A�CTAT5�� ����e"�USER��@�O�BT�@�CksT�C�T4�T5�T6�T�7�T8�Q*�NDO_CFG ,9�Xt�s�*�PD-QgY��None� *�^P_INF�O 1-�e`��0%�O,o�xo[o >oo�oto�o�o�o�o �o!EW:{�b��QOFFSET' 09�a�PC ��XO����/�&� 8�e�\�n��r����� ȏ�����+�"�4�F� ���ϒ�����
��ڟ��xUFRAME � PD�V�QRTOL_ABRT����s�ENB��G�RP 11�Ɋ�?Cz  A�u�s� �Qs���������ͯ߯���x�U?��Q.�MSK  B�a.�mN��%	i�%b����k�VCMR[�2�7�{#�R@	��Pfr1: S�C130EF2 Q*ݿ�PD�����T�&��5R@�Q?���@�p��ȇ� ɟ5�?�IH`�@rϟ�ı����8�屢A�RB���RB? B����RA #ի�Dߋ�h�7ߌ�w� �ߛ��߿���
�a��� @�+�=�v�)ߚ��ISIONTMOiU�B��U�����R8SﳸS�� j� F�R:\��\�PA\��� �� M�C�LOG�  � UD1�EX�5�RA' B@ ��x�I�r����I����PC �� n6  ��q�IFu�%��`���Z�  =����PD	 J�*�TR�AIN_���ǐ  dPp	�栲9�}(c��W� ������.�2@Rdv���_\�RE��:b�ʲ��/LEXE��;�{�Q�1-e��VMPHKAS/P�U�S����RTD_FIL�TER 2<�{ Ԓ��,�{/�/�/ �/�/�/�/�/??�� i/N?`?r?�?�?�?�?��?�?�?��SHIF�T�1=�{
 <��q�JODU)OOO�O _OqO�O�O�O�O�O�O _<__%_r_I_[_�_�_	LIVE/�SNAPesvs�fliv.�_���� �pU�P�Rmenu�_�_�_Woio�@b	E��>IO�EM�O��?�� ��$�WAITDINE#ND��+��dO?�"���g���oS�iTI]M@���<|G�o ^}�o�{az/azN�hRELE%!@��dx�����a_ACT�Pp�K�E�� @d��ko���E�RDIS��PA��`V_AXS-R�p2Ab������Vp_IR  +&�� 	��)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ��������XVR�aB~��$ZABCp;1C� ,N f�2ϵ�ZIP��D�e������ύ��MPCF_G 1Eٍ0J��=��S�qFىX�`# �c�܋߆�<90 ��߻�S�|��ߠ�?� }������S��$�z��8���� � ����������
�4�M����G��JÛ�YL�INDK!Hً �Є� ,(  *��������������� ��);M�� p���{���  U6��lS��w�����Y�29Iه]� �)�#/ 3,���\/G/�/��/��/���!A�c�S�PHERE 2Ju��*?z�/<?#? `?��/�?�?$�?k? Q?O�?&OO?\OnO �?�?�OO�O�O�O�O`EO"_4_F_M�ZZ/� ǘf