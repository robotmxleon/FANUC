��   ��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����BIN_CFG�_TX 	$E�NTRIES  $Q0FP?UNG1F1O2F�2OPz ?CNE�TG  �DHC�P_CTRL. � 0 7 AB�LE? $IPU�S�RETRAT��$SETHO�ST� �DN�SS* 8�D��FACE_NU�M? $DBG_�LEVEL�OM�_NAM� !����FT� =@� LOG_8	,�CMO>$DN�LD_FILTE�R�SUBDIRCAPC � �8 .. 4� H{ADDRTYP�=H NGTH��f��z +LSq� D $RO�BOTIG �PE�ER�� MASKn�MRU~OMG�DEV����RC�M+� 7�$ /�QSIZνTIMR� TA�TUS_/!?MA�ILSERV �$PLAN� <�$LIN<$C�LU��<$TOޥP$CCw&FR\w&YJECZ!8%�ENB � ALkAR!B�TP,Թ#,V8 S��$�VAR�)M�ONx�&��&APPL�&�PA� �%��'PO�R�7#_�!�"AL�ERTw&G2URL� }83ATT�AC�_0ERR_oTHRO33USt9&!u8� CH- A%�4wMAX?WS_Z1w��1MOD��1I� $�2M }(�1PWD  } cLA�r0�ND�1�TRY�6DELA�C�0%'�1ERSI���1/'RO ICL�K=HM� /'� XM�L+ �#SGFRM�33T� /!OU33P�ING_�COP��!�F3�A/'DUM�MY1�G2?���RDM*� $gDIS�!SM l5�M!n"Y%/7�ICC�%� �FVRe0GUP� _wDLVSPAR�O�SN
#	3 q_)R/!_WI�CTZ_INDE�3θPOFF� ~UR��YD��Sk  ?
 t 8!]P'MON� cD�bHOU3#EAf.axf.a%fLOCA� �A#$N10H_H-E���@I�/ }3 $ARP&&��_IPF�W_� O�F�PQFApQD0�VHO_� oINFOncEL�G P����0WOR�1$A7CCE� LV5[:02�ICE�'p��@�$�c  ����Fq��
��
�;p&PS�ADw�# ��WqIX0A�LCUq' dx
�
��F����op�r�uw�$� 2�{ "��Qr�}�p�� ğ}��!Mq5����$�� _FLTR  \cy�p ���������I�$�}2�I��bSHyPD 1}�y  P1�珴t֏��7��� [���B���f���ٟ ������!��E��i� ,�>���b�ï��篪� �ί�A��e�(��� L���p����ҿ�ʿ +��O��[�6τϩ� l��ϐ��ϴ����9� ���o�2ߓ�V߷�z� �ߞ߰����5���Y� �}�@�v���������M�z _L3A1�b�x!1.6�0����5�1F���2�55.~�=�����u4�2;�M���a�s�������3��M�* ��������4+M��  Qcu���5�M�@������6�M��ASew����$RC�`G �MA� MA���Ѐ�v� OQ� ���<-/ b/t/G/�/�/�/�/�/�/��P�/"?4?F?? j?|?�?�?_?�?�?�?��?��u2OLO��?wO�O�O�O��}�iRConnec�t: irc�D//alerts�O �O__*_�EqOV_h_�z_�_�_�_���sP�"��d���_�_�_ o!o3oEoWoio{o�o�o�o�o��$E_�o��(�oiO:L^pR����(�$"��r&J�u�q��� D�M���$SM&��ŋ��%1�D���I���8�q��\��� L�qN�q
!	��~��珿�p������ #��US?TOM 
�}����#  ���T�CPIP�r�}�$H%�TEL���u !� �H!T��R����rj3/_tpd�� (�ׁ?!KCL�����׏��v!CRT����W�"ߔ!OCONSX���őOsmon]�ߔ