��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A   �����
�WVAMP_�T   �$X1  $kX2AY@@/�FC5  �$2ENBA $�DT  / _�R2 d EN�ABLEDnSC�HD_NUMA �xCFG5�� $GROU�P�$z ACCE�L@�G$MA?X_FREQ�2 �L�DWEL�D�EBUG�PRE;WSOUT��PULSEAS�HIFt 7TYP�4$USE_A�EF} 4$GD=O�  f0� r?�NpW�EAVE_TSK� �V�_GP��SUPPORT�_CFnCNVT_DONE p �}k}GRP #2r�� _� ��$� TIME1�o$2'EXT�� (1#&(MODE�_SW�CO3 S�WIT � C/ P�HAX6  4 m� ECC$��TERMNnP�EAKno!AL ? \ � �!�I�$�!N_=VSTAR�#!�r"��"�%�C�YCL42 
���/ � Tv"b �$CUR_RELq_� �!3WPR5� � 
$CE�N� _RI3RA�DIU�XI�z ] ZIMU�Ti!$ELEV�ATIONg5� N��CONTINU�Oe2q �MEXAC=PE�S�6 � H~ �UEN�CYA�ITUD<4�2RIGHC�2�LEBL_ANG�1 �OTF_�� 	�  1$3A�bET���n3C!$O;RGjHFBKjH���P��C��DLD%W�HR�E�_�3�B �C��D�B�C�@�D�A�CCHG�G	Q�F	Q8�F	Q�FINC�G=Q �F=Q�F=Q�F�AVCPYC� _T�\#�Y�~P#�@SY��H)@�UPD"0n��$$CLASS  ����Q���8 �P�PVERS��1�W  ����QIRTU�AL�_�Q0 2~�X�  ��{?��@�  Ha Dae�TWoio{o�o�o�`)dN 2 3k� Hf��uHe@O�Hi�oNc)a� � e� E`���`9t12  �z����=�����4s ����jpYq��w�r��1��x at��ujp`��i.�5t8q�q2�b�t���
�9x��������̏ҏ���Sb�)a�  23k
=TDaSI�8�� �����0h�?m�'����l�D��� ��Ca��l����k���� �2�D�V�h�z��l�FIGURE 8��o�v�Hal� f��������M�(� H��󈯎�����Ŀֿ~�TCIR1��Pd�}�0�~�h�0z�D�Z�l���0�v� ��~����� ��$ߪjN� Hp��4q�Ȓ���@��ʖD�M` g����������	���-�?�Q�c�u�`�� �q� �5)�ᐟN`���ᬟ ����˟���M�_�q�������������k�Triangle��z�h߾�M�� Ɵ�ύ�����0�/ L� &��g�n�� �	//-/?/Q/c/u/ �}DVhz��/�/ ��9?K?]?o?�?�?�?�?�?����� O �h��O2ODOVOhOzO �O�O�O�O�O�O�O
_ _.[�?._O"O�_�_ �_�_�_�_�_oo&o�8oJo\ono�mSCH�EXTENB  �=��ctSTAT�E 2�k �|o�o�o �gWPR 7�6�L}D��-�_OTF 	8��@)0�q�q����v)��uAȫs�u@�  <#�
�?�����mu_GP 2w| ���d� v����я㏡+