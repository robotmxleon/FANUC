��   F��A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A #  �����#�AMON_D�O_T   �$PORT_�TYPE  �@NUMJ/SG�NL7 L�$MIN_RAN}GI$MAXr�NOo ALxp V��~ �COUNT>J �AWE08 �� $AWn0ENBJ $�|G1LY_TIV�$WRN_ALM�STP�
�E��C�.�WT�C�
J�AFT_�CHGxAVRG�_INT��{SgAVE�YP1?ER_REG�Tw$WA� SIG�� OP��V/OLTS�����AMP�&AEx �#E_VL� �&D'>% I*f$� _�ANL�  �p 
$US0 S�_CMD � PRIORITY�"�UPPER� $�LOW�$�#$FgDBK�"�RAv ~�!SQ_AVG�#n�#SD_� CE� r� O��$ �� � LIN�!$A�RC_ENABL��!� 0DETEC��!< ELD_SP~�$PD_UNI���!92DIS�"�I�D IM�#��  v1WFt2���CF�" � �$PS_MANU�F �2OD�EL�5PROCEySN0�0WFEEW0�ESC�2�2_FI�#1�1�1�7T _AOT�"�2I�6D�7DC`1�6L �"{2 � �CNV� 7   $EQ�zxvODOU� A<CkTBd� $?C? 2 �?@�DD   , �� MM�!�$D� ��!2� $F� �B�4NuV7	JBSEL10�_NOJDATA�_s@�@ {"W�PpG
{M
�FWP�7 L@�L
 ��WIR_CLP4 L@AS�BU8  H $(4��R�4�YPREF� �U;A�_ECU��  �JB~ �S  � $BPEEPf#�}!SCH7 � �!��`�1e�#dPK*jFRE�Q.gULSwbSP�0fg2y�!hyb�*g�F�AI6 �ZCoVG}�hp  dD�e�e�`�	�a��d�BVB�aZERO8y}uSLO]R�`NT�!P�cO	U\93|�L FORMA0�NAra�0J3	�� D�cQWUXW�EIOEX7'4 �A�WfxccmpS_91INp�� :1�U�p� FA1UG"t0LO�0�q�P�!�G��R<�A<Dp;�STIC�@�p�ROBOT�AD�Y�rERRO�S�E��`S��p�!T�R��$S�CHDO�G_�@%��0_AC�TIV���I�Cʯ01�2�q�OT�F7 � $ 
��P��x�nfpNCi0�c;�f 0�*d;�*g0�7f;�7i 0�Fd;�Fg~�Td��Tf�UP�@�B�sPCR�7�� WSTK��� =�Hr ՒƁ %��00��2�X���0�A~�3KIPTH�E91�S;������PIKEf���0�0�WWV�2t�E_HaO;0�0��PHK-18���� RMT����SPTL�0p�$�Hz��SW��pd�$BBg1_ONL4�$B�2pf�bgF�WF�1e2_R��0zE"�!� _W;6�A?ND1OFF���!�ND2g�3g�R�Sp� �A� �SEPM�? | $�0�@ g��e��*f��7b���Ff�TfADAPTz� G�CSENS��c��!ݒ��8 � 0?,2���"��$ �1b�!c�7cc�Fa|� Tac�^��'y��&l��&*�!4�&5�&6�"8��W�@�2 HOU�!h�o � �SE�0 �g4�Q�T<��6��'��46�q56�0� ?%$CURR7(�^�"HEATzPe@ �!燰"j���i�p��GAP�#Ti�XPY0���EHP��@��pDS��@�!GP�0S�!�$���$GO� RI����AM�#/"�#M䩰jAN3O�BEFB ;�LHV1[5j�� 43;1 `H�V�PA�H�r���3��F1�� _P�/�SR 7 �+ 	� RSB�$�� 0G�m�b�O�J���O��DU�IW�A�XQl�2C,1L�"D�����?3���8 � 4�@P֋q]ִSG�ʦ�~�;A8�8  $ $�@�CL�$ć�s	۔��8 $ ;o2� �"�ql�0�q��� 	PK�P�� 
��*���q�BPa��b�@4�5�6:2K�3���&��FW�q�B��ALAR���2��2@�����
�3�Q_R}��
�.4�4�F�+�PW,���_ @ĸ�Ӕ]���� ���Qbwm��t���QDI�c�j��~pus��R�SIZ���BGOAR���1]E7�]�\�h"0h"��ķ�$VEN�D��I��DEVI�C��0D����MA5J��V�#IN�(�$�uI"�vMA��p�FI�0�BW����� p $��X��h ⡡��F̀OR_R���C�^1D4TO_l��O5_R�pRS<�f'�OS�9�BUP� #N�:��0 �`�=� �6��6��9�PURG��RKtS�TFR�p&���A ��.E�.E�AED��P$-��M%�fMT�����eEM7��Q�5��� Z$�22�9�P駇��K��p�QADJ�T��NsEXT��r_LE�c"��P��X��M����aA��_�#IV���1H�q�2�eFL������P��:����0�8� ̀�;�WT[�CY��� ���q�  �	`��`( ~�bTOTAL_�Qȑc���VI�p�WWARo��U��A*�P1Y&1b�uKG����'" A}�#N�p { �SCFG�1wz�LOO�B:��P�Q�S!@���GLOB�P�⣠ܽ ��NOT��$b0QI4�*��AVh�Y��$��������e���W_SHFL�W�X�fkrI�$�q �e�RY	��оP��%�ʀLIMS`�i�@��c7�UIF�e�A�PCOUPL�R @ �p�q���[ �qUR�`N��<�MMYm �u0̼u�  ����US�TOk�   � x�0 �qp` �
  ��SEMG�g��1! ,��MGX�Ag���NOzPR ���wa�"� ,/���Ȣ=6Ƞ��3T� )�RT���p�0=����AHER� A�������'"݈{�� �����@���Q�L�� )BD ��2C���7B<�^i3_FIL@�W��7BUG_3SM ���ñF_F����q�, �_4N SV@БTC�P��=Ҕ�DIO��������.a�TM�C��PA�Pq��q�w�x��q�_DYN�V�2Wԣ����KE�YV�GQׂ��F`��?�/B�{�_C��R�TOU���������CAL�Q0�`�� TIp1�P_y�R�T���@��A?2 ��$$CLASS  �������� �-�S�B���  ����IRTUx�����AWAOY1h��[�$�
��K���n�2�f��[�[���g�
�?�������g������� ����(�:�L�^�ppςϑ�l�EXEu� `���������Ͽ�*� <�N�`�r߄ߖߨߺ�\��r@S Rw��� :����#�5�G�Y�k� }���������������l�NLG 2Mx� �����?�ˑ<1�6�`��e��� pp`����{` 2:��)�Ge�neral Pu�rpose��MIG (Vol/ts, 0)���� ����
AWMG�ENL.VR�A*EGLMG19��g�`������ ��'���������������CNV� 2	x��[������ 4aPzUh�� ���//�=/O/ ./s/�/\�/�/b/�/ �/�/?'??K?]?<? �?�?r?�?��E�/�? O�?2ODO#OhOzOYO �O�O�O�O�O�O
__ �?@_R_�Ov_�_g_�_ �_�_�_�_�_o�_(o No�?ro-_�o�o3o�o �o�o�o8J) nM_�{o��� ��� �F�%�j�|� [�������֏�go�� �0�B�!�f�E�W��� {���ҟ������,� >��b�t�������� ί௿�����:�L� +�p����O���ʿU� � �߿$�6��Z�l� KϐϢρ����ϯ��� ߵ�2�D�#�h�z�Y� ��}ߏ��߳���
��NVWP 2|	:i\>�T 
��b��t���USTOM� 2|l  A��������h�	h�d"���DEFSCoH R|�Q��<�b�@Default Schg� ��n��������� ��K"4�Xj �������
)��FBKLOG1 �@��T�῀ � Ugy��12�=O����5L�G_CNT  �����)�IOEX k2�����A ��+C�]$@�������!�
Weld� Spee%��IPM  d$�/�/��/�/??(?:?��O_TF 2��A?��?�?�?�?�?C8=7�����@����?�K)�PCR 2���pI�BH�?��B�C!�FK<D7�*��>��?�ffAZ �A�"��OFM"@�����/�O@O"@.�����WOELGG��k%*_�F�0�2345678901JRUK%4_y_�_ĝ_HIȩ_7]�OOS�RAM2��IB�$��_oCRGSEL� R<�Q� �	Process# 1oSf2�_ojU3i�o4i�o�5�-mlXS���o7���kn8i'l"@>��� �_);E�s-B� �W�%�Voltage���qsfc%Dw<|!@]y�h����aWire� f�  s�$	 � hc%[&t/�oDS� l*�<�N�`�r����� ����̏ޏ����&��]+zvd"����  ?�#��E�Z"!���a��^/�� ���V���a�aɒCurrent�Amp�=���l �eu���Q�c�u����� ����ϯ����)� ;�M��W���a������ ��	q��)q��Iq��R� ͹ϧg�a�aA��b-� ��-�	q-�)q-�VE!���\e�	q?���*�Z�%�������ϻ������PDRuS3 R\zH��jq��C�U�g�����gߩ� ��u߇ߙ������� ��]�o�)�;�M���� �����#������ k�}�7�I�[������� ����1C��I ��Wi���� ��?Q/� �����//)/ ;/M+�U/g){/�/�/�M/�/?cS2�S^=�R��b�S2UPYp�^=�=�o?��33H1>E0=L�S�>I0h!�@"�@�#�@$�1t9�g�$q�#?�v�#>�8�8�CWIRE 2�&M<�?�?h�>��3�>�G(=��J*�ESCFG �G�A��Y��OO��E7])COUPL*�0=k
0�vk B`�D�^�L�[�OZW�O��G_�OP_G_Y\�HN�B  ��Ec&FUSTOM  =k�
8ƙy�O&EEMG?OFF !=kS���)BPCR �"�_��@���zqC {sUūMJo�\zt�f_oeo��
Cl�q¨1