��   v1�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����UI_CONF�IG_T  � E$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]5�ODE�
6CWFOCA �7C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"�%�!BA�!j ��!�BG�#�!hINS�R$IO}7P}M�X_PKT?$IHELP� {ME�#BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�<ST]Yf2$Iv!_Gv!k FKE�E ��8C &USTO}M0 t @;AR$@PIDDbB�ChD*PAG� ?�^DEVICEބISCREuEF���}GN�@$F7LAG�@ KB��1  h 	$P�WD_ACCES � =EFB�S:1~�%)$LABE� O$Tz j�@��32R�	&U�SRVI 1  < `'R*'R�n(QPRI�m� �t1�PTRIP�"m��$$CLA�@ �����Q��R2��R�P\ SI��W�  �׸QIRTs1�_�P�'2 L17�L1�A�R	 ,���?���a�P($bda����`�� Ao��
� ��'/SOF{TPb@/GEN�1�?CURRENT�=>�A,18,1 lo�o�o�o�o �o�o,95,2�o?Q�cu �(5 �`w�����)q9�G�Y�k�}�� ��s�oˏݏ����>��E,381�oN� `�r�����Q������ ӟ���	���-�?�Q� c�u��������ϯ� ����)�;�M�_�q������aTPTX��&���˿`� s����$/�softpart�/genlink�?help=/m�d/tpmenu.dg��2�D�V�h� !��Ϟϰ�������u� 
��.�@�R�d���u� �߬߾������߃���*�<�N�`�r������Q[f=bOb�� ($��������������Qa:�<cI�<c:�8����zc��RBa��>a�����  ��	����%����`�[`^��W`  ��� ���SQB 1~�XR \���_�� REG VED��FX�wholemo�d.html	si�ngl}dou�b�trip��brows �t�Y��C Ugy��C-g�ydev.s�lh/� 1,	t0/ �/��/�/�/m/��/�/�/�/?8?� �PP?b?t?�?�?�? �?�?�?�?�6�@M?"O 4OOXOjO|OKE;	3? -?�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_�oo3o EoWoio{o�o�o�o�o �o�o�o/AS ewE?����� ��0�B�T�OOx��� Y�k���ҏ�O�O�� �'�9�b�]�o����� ����ɟ�����:� 5�G�og�a������� ůׯ�����1�C� U�g�y���������ӿ �� �2�D�V�h�z� �Ϟϰϫ����ϵ��� �.����ݿv�q߃� �߾߹�������� %�N�I�[�m���� q���������!�3� E�W�i�{��������� ������/��j |������� �0B#x� A�S�9����/ /'/9/b/]/o/�/�/ �/�/�/�/�/�/��? ?G?Y?k?}?�?�?�? �?�?�?�?OO1OCO UOgOyO�OY�O�O�O �O_ _2_D_V_h_c��_�_m__�_�_�Z��$UI_TOPMENU 1�P�aR 
�da�A)*d?efault�O�M�*level�0 *�K	 �Ho60�o/o�o�btpio[23]-8tpst[1�h��o�o�oko}o(=h�58E01_l.�png</6me�nu5^yUp�q13^zr]z}t4�{l)q����
��.�@� R��B�{�������Ï�Տd�prim=��qpage,1422,1܏�'�9� K�]�h���������ɟ�۟j���class,5��+�=�O�4a�l���13h������¯ԯ�m���53�"�4�F�X�j�m���8�����ɿۿ �l��#�5�G�Y�k��I`a.o��Rm��`+q������fty�m<�o�amf[0�o��}	�c[164�gf�59�h+q�ߣ�yx2��}�ҙz��w ]{��s����n��� �����������"� 4���X�j�|�������A���2����/ A���w���� N`�� $6H��	�1\������M���ainedi��//)/;/M/�H�config�=single&>��wintp��X/ �/�/�/�/�Ja���/ ?Se?%��E?W?i? |?�?�?�?�?1?�?�? OO/OAOSOeOwO� �O�O�O�O�O__M� >_P_b_t_�_�_'_�_ �_�_�_oo�_(oLo ^opo�o�o�o5o�o�o �o $�oHZl ~��1���� � �2��V�h�z��� ����?�ԏ���
��.��N��d��������ϑO��5�s�̟�'�ٗuݤ��� ������3��ڂ�����̩6ٯu7�F�X�1�C� U�g�y�ď������ӿ ������-�?�Q�c�(uχ�f"\1k�� ������	��-�?�Q� c�u߇�߽߫����� ����Z�M�_�q����$�6�6������`����d$�74$� U�g�y������,C����5	TPTX[2c096��4��246�0������18"P4F��0�25�`�1��i���tvԡ�����0�1����C:l$tre�eviewy#�3�C�&dual=o��81,26,4 $�����//// A/S/e/��/�/�/�/��/�/&�;x�53 ��E�O?a?s?~/�? �?�?�?�?�?�?O'O�9OKO]OoO�/?:�1�%?�2���O�O�O �6�O.�edit ��O�OT_f_x_'�w 5�1_CS�_�_�_o�� o4o�<o�Uo!{o �o�o�o�o�o�ogo /ASew�� ������"�4� F�Oj�|�������ď S������0�B�я T�x���������ҟa� ����,�>�P�ߟt� ��������ί]��� �(�:�L�^����� ����ʿܿk� ��$� 6�H�Z�	oo��?o�� �������� �1� C�U���aߋߝ߰��� ������	��@�R�d� v������������ ��*���N�`�r��� ����7������� &8��\n��� �E���"4 �Xj|���� S��//0/B/� f/x/�/�/�/�/oρ� �/��?���=?O?a? s?�?�?�?�?)?�?�? OO(O9OKO]OoO1� �O�O�O�O�O __]/ 6_H_Z_l_~_�__�_ �_�_�_�_o�_2oDo Vohozo�o�o-o�o�o �o�o
�o@Rd v��)���� ��*��N�`�r��� ����7�̏ޏ���� &��/�/\�?���?�O ����ǟٟ����!� ��-�W�i�{������� ïկ�O��0�B�T� f���x�������ҿ� �����,�>�P�b�t� ϘϪϼ������ρ� �(�:�L�^�p߂�� �߸������� ��$� 6�H�Z�l�~���� �����������2�D��V�h�z���:�H�*default���j�*level�8�M��	�� �tpst[1�]	KyPtpio[23R6H�uP����m�enu7_l.pkng��13�	B5
��41u6�
�w��� ����//+/=/ O/�s/�/�/�/�/�/��/n"prim=��page,74,1�/?-???Q?c?�n"�&class,13h?�?�?�?�?�?u?�25�?"O4OFOXOjOm#|<O�O�O`�O�O�O�/218?�)_;_M___q_|O�26�x_�_�_�_�_�_���$UI_USERVIEW 1J��J�R 
��EDIT�,Weld DA�TA s�dou�blej���_�medit1eo�oФo�o�okj�&95 P�o,>�o�o�t���p�0cST�ATUS,POS@ftripMo_oqo@�,�>�P�b��Yy�2m�����ÏՏx�33_��1�C��P� y�t������˟ݟ� ���%�7�I�[�m�� ������ǯٯ����� 
�|�E�W�i�{���0� ��ÿտ���Ϯ�/� A�S�e�w�"��ϖϨ� �������+���O� a�s߅ߗ�:߻����� ���ϸ�"�4��X� �������l����� �#�5���Y�k�}��� ��L������D� 1CU��y��� ��v�	-? ��L^p���� ���/)/;/M/_/ /�/�/�/�/�/v�/ �/�/n/ ?I?[?m?? �?4?�?�?�?�?�?�? !O3OEOWOiO?vO�O �OO�O�O�O__�O A_S_e_w_�_�_>_�_ �_�_�_o�R