��   ��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����BIN_CFG�_TX 	$E�NTRIES  $Q0FP?UNG1F1O2F�2OPz ?CNE�TG���DHC�P_CTRL. � 0 7 AB�LE? $IPU�S�RETRAT��$SETHOsST��NSS*� 8�D�FA�CE_NUM? �$DBG_LEV�EL�OM_NAmM� !� FT�� @� LOG�_8	,CMO>�$DNLD_FI�LTER�SUB?DIRCAPC���8 . 4� H�{ADDRTY�P�H NGTH���V�z +L�Sq D $?ROBOTIG ��PEER�� MA�SK�MRU~O�MGDEV��R�CM+� �7$ /�QSI�Z�TIMR� T�ATUS_/!?MAILSERV� $PLAN� �<$LIN<$�CLU��<$T�O�P$CCw&F�Rw&YJECZ!�8%ENB � A�LAR!B�TP�,�#,V8 S���$VAR�)M�O�N�&��&APPL��&PA� �%��'P�OR�7#_�!�"A�LERTw&G2UR�L }83AT�TAC�_0ERR�_THRO33US0t9&!u8� CH- A%�4MAX?WS_�Z1��1MOD4��1I� $�2M �(�1PWD  �} LA�r0�ND�1TRY�6DEL�AC�0%'�1ERS�I��1/'RO IC�LK=HM� /'� X�ML+ �#SGFReM33T� /!OU33�PING_�CO�P�!�F3�A/'DU/MMY1�G2? �DM*  �$DIS��SM l5�M!�n"%/7�ICC�%H� FVRe0GUP� �_DLVSPAR��QN
#	3 �_)R/!_WI�CT?Z_INDE�3�PgOFF� ~UR�Y�D��Sk  
� t 8!]PMO�N� cD�bHOU3#EAf.af.a�%fLOCA� A#{$N10H_HE�K��@I�/ 3 �$ARP&&�_7IPF�W_ O2�F�PQFAQD0��VHO_� IN�FOncEL� �P���0W�OR�1$ACC�E� LV5[02��ICE�'p� ��$�c  ��)�Fq��
��
;p&PyS�ADw# k��WqIX0ALC�Uq' dx
���F�����op�r�u�]$� 2�{�@ ��Qr�}�p�� �}��!Mq5����$� _?FLTR  cy�pW �������!�I�$�}2I��b{SHyPD 1�y  P1�珴t֏��7���[�� �B���f���ٟ���� ��!��E��i�,�>� ��b�ï��篪��ί �A��e�(���L��� p����ҿ�ʿ+�� O��[�6τϩ�l��� ���ϴ����9���� o�2ߓ�V߷�z��ߞ� �����5���Y��}� @�v��������M��z _L3A1b�x/!1.6�0����5�1F���2551.~�=���ܼu4�2;�M���a�s�������3��M�* ��������4+M�� Qcu���5�M�������6M���ASew���$R�C�`G ��� ˷��Ѐ�v� Q� ���<-/b/t/ G/�/�/�/�/�/�/��P�/"?4?F??j?|?��?�?_?�?�?�?� �?��u2OLO�?wO��O�O�O��}iR�Connect:� irc�D//alerts�O�O_ _*_�EqOV_h_z_�_(�_�_���sP�"��d���_�_�_o!o 3oEoWoio{o�o�o�oD�o��$E_�o��(�o�iO:L^p����(�$"�r&Jd�u�q��� DM����$SM��	ŋ��%1�D���I���8�q�\���$ L�qN�q
!	�~���珿�p������ #��USTOOM 
�}����#  ���TCP+IP�r�}$H%.�TEL��u !=� �H!T�R�����rj3_t�pd�� (�ׁ!KCL����׏��>�v!CRT����W�"ߔ!CO�NSX���ősmon]�ߔ