��   v1�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����UI_CONF�IG_T  � E$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]5�ODE�
6CWFOCA �7C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"�%�!BA�!j ��!�BG�#�!hINS�R$IO}7P}M�X_PKT?$IHELP� {ME�#BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�<ST]Yf2$Iv!_Gv!k FKE�E ��8C�&USTO}M0 t @;AR$@PIDDbB�ChD*PAG� ?�^DEVICEބISCREuEF���}GN�@$F7LAG�@�KB��1  h 	$P�WD_ACCES � =EFB�S:1~�%)$LABE� O$Tz j�@��32R�	�CUSR�VI 1  < �`'R*'R�(QPRI�m� t1�P�TRIP�"m�$�$CLA�@ �����Q��R��R̜P\ SI��W  �׸QIRTs1�_�P'2 �L17�L1A��R	_ ,��?2���a�P$bd�ab��`��  ����
 ���'/SOFT�Pb@/GEN�1?�CURRENT=|>�A,18,1lo��o�o�o�o �o�o,95,2�o?QcNu �(5�` w�����)q9�G�Y�k�}��� �s�oˏݏ������E,381�oN�`� r�����Q������ӟ ���	���-�?�Q�c� u��������ϯ�� ���)�;�M�_�q������aTPT�X��&���˿`� s����$/s�oftpart/�genlink?�help=/md�/tpmenu.dg��2�D�V�h�!� �Ϟϰ�������u�
� �.�@�R�d���uߚ� �߾������߃��*�`<�N�`�r�����Q�[f=bOb�� ($��������������Qa:�<cI�<c:�8����zc��\a���>e��  ���	������Ģ�`�[`^�W`  ���� ���SQB 1�XR� \��_��� REG V�ED��FXwh�olemod.h�tml	singl�}doub��trip�brows�t�Y ��CUgy���C-gydev.s�l/� 1,	t0/�/� �/�/�/m/�/�/�/8�/?8?� �PP? b?t?�?�?�?�?�?�?�?�6 @L?!O3OO WOiO{OJF;	3?-?�O �O�O�O�O	__-_?_ Q_c_u_�_�_�_�_�_ �_�_�oo3oEoWo io{o�o�o�o�o�o�o �o/ASew E?������� 0�B�T�OOx���Y�k� ��ҏ�O�O���'� 9�b�]�o��������� ɟ�����:�5�G� og�a�������ůׯ �����1�C�U�g� y���������ӿ��  �2�D�V�h�zόϞ� �ϫ����ϵ����.� ���ݿv�q߃ߕ߾� ���������%�N� I�[�m����q��� �������!�3�E�W� i�{������������� ��/��j|� ������� 0B#x�A�S� 9����//'/ 9/b/]/o/�/�/�/�/ �/�/�/�/��??G? Y?k?}?�?�?�?�?�? �?�?OO1OCOUOgO yO�OY�O�O�O�O_  _2_D_V_h_c�_�_�m__�_�_�Z�$U�I_TOPMEN�U 1�Pa�R 
d�a�A)*def�ault�O�M�*level0 =*�K	 Ho60�o/o�o�btpi�o[23]-8tpst[1�h�o�o�oko}o(=h58�E01_l.pn�g</6menu15^yUp�q13^zr�]z}t4�{l)q�� ��
��.�@�R��B �{�������ÏՏd��prim=�qp�age,1422,1܏�'�9�K�]� h���������ɟ۟j����class,5��+�=�O�a�l���13h�����¯hԯ�m���53�@"�4�F�X�j�m���8�����ɿۿ�l���#�5�G�Y�kϖI `a.o��Rm��+q������fty�m�o�aOmf[0�o��	Пc[164�gf�5�9�h+q�ߣ�yx2 ��}�ҙz��w]{� �s����n����� ��������"�4��� X�j�|�������A���2����/A�� �w����N` �� $6H��	�1\�����M����ainedi���//)/;/M/H��config=s�ingle&��wintp��X/�/�/ �/�/�Ja���/?Se ?%��E?W?i?|?�? �?�?�?1?�?�?OO /OAOSOeOwO��O�O �O�O�O__M�>_P_ b_t_�_�_'_�_�_�_ �_oo�_(oLo^opo �o�o�o5o�o�o�o  $�oHZl~� �1����� � 2��V�h�z������� ?�ԏ���
��.��N��d��������ϑO��5�s�̟�'�ٗuݤ��� �����3��ڂ�����̩6ٯu7�F�X�1�C�U�g� y�ď������ӿ��� ���-�?�Q�c�uχ�
f"\1k������ ��	��-�?�Q�c�u� ��߽߫�������� �Z�M�_�q���$�6�6����������d$�74$�U�g��y������,C���5	�TPTX[2096��4��246�������18"4F��0�25��1��i���tvԡ��$��0�1����C:l$treev�iewy#�3C�&�dual=o�8?1,26,4$� ����////A/S/ e/��/�/�/�/�/�/2&�;x�53�� E�O?a?s?~/�?�?�? �?�?�?�?O'O9OKO ]OoO�/?:�1%?��2���O�O�O �6<�O.�edit��O �OT_f_x_'�w5�1_ CS�_�_�_o��o4o �<o�Uo!{o�o�o �o�o�o�ogo/ ASew���� ����"�4�F�O j�|�������ďS�� ����0�B�яT�x� ��������ҟa���� �,�>�P�ߟt����� ����ί]����(� :�L�^��������� ʿܿk� ��$�6�H� Z�	oo��?o��� ������� �1�C�U� ��aߋߝ߰������� ��	��@�R�d�v�� ������������� *���N�`�r������� 7�������&8 ��\n����E ���"4�X j|����S� �//0/B/�f/x/ �/�/�/�/oρ��/�� ?���=?O?a?s?�? �?�?�?)?�?�?OO (O9OKO]OoO1�O�O �O�O�O __]/6_H_ Z_l_~_�__�_�_�_ �_�_o�_2oDoVoho zo�o�o-o�o�o�o�o 
�o@Rdv� �)������ *��N�`�r������� 7�̏ޏ����&��/ �/\�?���?�O���� ǟٟ����!���-� W�i�{�������ïկ �O��0�B�T�f��� x�������ҿ����� �,�>�P�b�t�Ϙ� �ϼ������ρ��(� :�L�^�p߂�ߦ߸� ������ ��$�6�H� Z�l�~�������� �������2�D�V�h��z���:�H�*de�fault��j�*level8��M��	�� tpst[1]	�KyPtpioG[23R6HuP�����men�u7_l.png���13�	5�
��41u6 �
�w����� ��//+/=/O/� s/�/�/�/�/�/�/n"�prim=�p�age,74,1��/?-???Q?c?n"��&class,13h?�?�?�?�?�?u?�25�?"O4OFOXOjOm#|<O�O�O�O�O�O�/218?)_;_ M___q_|O�26x_�_�_�_�_�_��$U�I_USERVI�EW 1J�J��R 
��EDIT,W�eld DATA� s�doubl�ej���_�medit1eo�o�o�o4�okj�&95P�o ,>�o�ot���p�0cSTAT�US,POS@ftripMo_oqo�,�P>�P�b��Yy2m�`����ÏՏx�33_ ��1�C��P�y�t� �����˟ݟ���� %�7�I�[�m������ ��ǯٯ�����
�|� E�W�i�{���0���ÿ տ���Ϯ�/�A�S� e�w�"��ϖϨ���� ����+���O�a�s� �ߗ�:߻�������� �ϸ�"�4��X��� �����l������#� 5���Y�k�}�����L� ������D�1C U��y����� v�	-?��L ^p������ �/)/;/M/_//�/ �/�/�/�/v�/�/�/ n/ ?I?[?m??�?4? �?�?�?�?�?�?!O3O EOWOiO?vO�O�OO �O�O�O__�OA_S_ e_w_�_�_>_�_�_�_ �_o�R