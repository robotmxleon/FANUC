��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����WVSCHD_�T   H �$FREQUEN�CY  $A�MPLITUDE�@DWELL_R�IGHTNLEF~]L_ANGLM�&EXT- 8� $ELEVA�TION@ZIM�UTH@CENT�ERX SMRAD�IUS@OG�$�$CLASS  �������z��� VERS���  ����IRTUAqL��' 2 ��� 
 ?��  @;=���BB�  :L^ p������.�  2)��1/ C/U/g/y/�/�/��'G  �	4�/�/ �!