��   K�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_���$$C�LASS  ������D��D�VERSION�  �VIRTUAL�-9LOOR qG��DD<x$p?������kn,  1 <DwX< y�����C�����	/��	Z�Zm//�/�_/�/�/�/$ ��/�/	?';�$MNeU>A\"�  <��4/d?��[=-/~�;�i� CI�?ܣ?�;DD@#����?�?{9@ 'v?@ CF�3O�?[O�= cO�OwO�O �O�O�O�O_�O_E_��;5NUM  ����� tUT�OOLC?\ 
xY?O�_Cj��GO �_	o�?o?o%o7oYo �omo�o�o1_�o�o�o �o;!CqWy �����sV�Q�V y�Wy