��  U��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A0  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ���AIO_CNV�w l� RAC��LO�MOD_T�YP@FIR�H�AL�>#IN_O�U�FAC� gINTERCEPf�BI�IZ@!LRM_RECO"w  � ALM�"�ENB���&ONܢ!� MDG/ �0 $DEBUCG1A�"d�$3A�O� ."��!_IF�� P $E/NABL@C#� �P dC#U5K�!M�A�B �"�
� O�G�f d��APCOUPLE, �  $�!PP=_D0CES0�!e8�1�!��R1> Q�� � $SOF�T�T_IDq2TOTAL_EQ� 3$�0�0NO�2U �SPI_INDE�]�5Xq2SCRE�EN_NAM� �e2SIGN�0�e?w;�0PK_FI�0	$THK�Y#GPANE�4 �� DUMMY1"dJD�!UE4RA��RG1R� � _$TIT1d  ��� �Dd�D� �Di@��D5�F6�F7�F8
�F9�G0�G�GPA�E�GhA�E�G1�G �F��G1�G2�B!SB�N_CF�!	 	8� !J� ; 
2L �A_CMNT�?$FLAGS]��CHE"� � EL�LSETUP �
� $HOMEm_ PR<0%�S�MACRO�RREPR�XD0D+�0���R{�T UTOB� U�0 }9DEVIC�CTI�0�� �013�`B�Se#VAL��#ISP_UNI�U`_DODf7{iFR_F�0K%D13���1c�C_WAxqda�jOFF_U0]N�DEL�hLF0pEaA�a7b??a��`$C?��PA#E�C#sATB�d�� oW_PL�0CH/7 <� PU�P��B
2ds�`QgdsD�UT�PHAgpS�F���WELD|H2/0 =Lc�7w7atAING�0�$�r�1�@D2�4%$�AS_LIN;tE��w�t_��2UCC�_AS
BFAIL��DSB"�FAL�0�AB�0�NR�DY��P�z$�YaN�Wq<��`DE6r ��`���+�����tSTK��+�;s7�;sNO�p��[�̈́r��U* Ȁ%�9 � ��  ��q`�G�C�G�+�U�S_FT�vpF�ǂG��SSF��PAUS����ON7xǓHO5U�ŕMI�0�0�ƔSEC�2�ry�i �rHEK0�v8vG#AP�+�	�I� � gGTH���D_I���T= �l���� �`�s9!̅����9!G��UN1���q���#MyO� �cE � �[M�c����RE�V�B7��!XI�� �R  �� OD�P-��dPM� %�;�/�"8�� F�q��
aX�0DfT p{ E RD_E%�~Iq$FSSB�&_$CHKB�pEde#AG� �p�  "
�$Ա� Vt:5���3�Mpa_EDu �� � C2��qS��`�vl �d$OP��0�2�a<�_OK<��Y�TP_C� <�pd�vU �PLAC��^}��p� xaCOM	M� �rD|ƒ��0�`��KO]B BIGA�LLOW� (tK�w�0VAR��xd!�1}!�BL�0S � ,K|a�r�PS�`�0M_O]|=՗�CCG�`=N�! �� ��_I_��� �0�� �B.��1S� ~�CC'BDD�!��I����0�@��84_ CCWp` OOL
��P'�M�M
�n�CHs$MEAdP�d`T�P�!���TRQ�a�CN���FS3��ir�!/0_F��( D�!��v CFfT X0�GRV0��MCqNGFLI���0UJ�p����!� SWIl��&"D�N�P�d��pM~� � �0EED��!��wPo��`�PJedV
�&$�p��1``�P��ELBOF� �=��=�p/0���3P�� ���cẐ�G� �>A0WARNM�`ju���wP��𼠤 CO�R-�8`FLTR^juTRAT Tlp�� $ACC�rT�B� ��r$OR1I�.&��RT�P�p\gMpCHG@I��E3�T{�1�I ̉ra�HK��� �����"�Q���HD(���a�2
BJ{PCT��3�4�5�U6�7�8�9�!����COfS�_rt���3�V�O�LLEC��"MULTI�b
2��A�
1c�O�0T_�R � 4� STY(2�R���).��pp�b�n� |A0@6Kb�Ib$���P�c���UTO=�cE�EXT!Y�
B�!�Q 2 
l��a0��Rpub����  �" ���Q����qc��~#!|��1Y�M�
�P8$  lT}R�� " Lqࠊ/��P��`AX$GJOB׍��W�';IGx# d��? %?78��3�p%���9_MOR��$ et��FN�
CNG&AF�TBA���6䱀JC��9��D@r��1CUR.KPa`/Ek��%��?��ttaoA4��XbJ��_R��|rEC�LJ�r�H�LJ��DA���I�����2G���]QCRfT&�C ��bG����HANC6$LG��iqda��N�*�Ya�Cᇁ�0|rf�R'L±�mTX���nSDB�WnSRA�SnSAZ��P�X��$  ' FCYT��e�_F��Pn�Re�M
P�QIkOh ������1��e����Cg���A���MP�a� ��HK�&AE�Up�p�Q�QI�'�  ]PI���CSXC��Zq( �xs��s��T�R�C�cPN����MG�IsGH"��aWIDR��$VT�P��9�E�F�PA cI�X�P,aQ�1u�CUS�T��U��)R"TI�T����%nAIOV����P_�L����* \q���OR��$!�q���-��OeP��jЅpIp�Q�u��J8�
��0�_�~}pPXWORK��=+�$SK0���nWADBT)PTRw�_ , �l@Ab��s�R0�ؠD��A:0�_C����=�+`H�PL�q��R�A�"��#�D��r�����BJ�b��9�����DB�Q2��-�r~qPR��ΰ�
x ct��. p�E�S�a� �LӉI/��-�( ��0���j� 1%��EsNE���� 2D��b��q	����3H�PC�  .$L��/$Ӄ�����gINE׶�q_D����ROS��E0"2`q��f0�p��PAZ�|tAsbETURN�����MRQ2UA@�C�RŐEWMwp��S�IGN�A&rlPA���W�`0$P�f1$P�P� 	2j���q����!��DQ��f������׶GO_AW;0���pvp��qajDCS'����CYx42O�1P�8�8���2��2��N�@��CtDۣDE�VIѐ 5 P7 $RBֳ���I�P.�i�I_B�Y�q���T�A9�H7NDG�6���x����b�DSBLr3�ͳ��aܢLe7 H �� ���TOFB̶�FE@Бg')��ۣ�f8��cDO�a�� MC9�@�"�`�sr�(��H�P�Wp�X�ܢSLAt4���9IINP!���� ж�ۡ�:D *�SPNp�#�@lƍ�1��W�I1��@J��E�q87�qW�N�NTV#��V n��SKI�STE^�`�b��pڥ�aJ_�Srjb_>���SAF��k���_SVBEX�CLU��po�D�pLX ��YH��%qΉ�I_V9`�bPPLYj���������_ML��L�VR�FY_D��M�IO�`  P�%`�b�Oe��LS�|b��%4}������aP�u���Y�AU NFzf�����)��#"�cD�4Ͱ� S��r�AF� CPX٣e�_� ;j��pTqA#���  ��SGN��<��<@3� P��c_�t�a���qd��rt��`UN>�����<@rD�p]�T`��`��%`����zrEF�p]I>�= @��F��\t6@OTS����|�������孂y Mr�N�IC>2K�GM A���iDAY�sLOCAD���D��5��o�EF pXI�%?j���~cO� �5�_RTRQU�@� D����0Q�p �EԠ��� �?K�%>`� ��GAMP*Pp��A�"�'; DB'��VDUtS�U��CABU�B`�NS9@ID�1WR$�Q!`�V[�V_#� ; ��DI@J$C� �/$VS�SE�#T �BDC�A� ���|�DBf�AE_�;VE�P�0SW!�!�@�x�3�� @�`�O�H�@PP <I	RwqDBB�p�=�!pU����t"BAS�рo'~P�Pn%[�d� B�	� ���RQDWf]%MS� �%AXC'<�;LIFEC���� ��	2N1EB5��D3EBCd@/Ź�Cq`ʡN�4q�6��3OVՐ%6HEh�DB'SUP�1��	2D�_�4j�H1_!C�5š
�7Z�:W�:qa�7�S��"BXZ�PʁEA+Y2HC��T�pސ��NM��zr0P�dgD `L��@HE�VXCSIZ?6k0��[��Nh�UFFI�0���C��������6ܭ�HMSWJEE �8��KEYIMAG�TM���S�A5���F���r��OCVI9E �qF 	�P�LQ�_��?� 	��&`KDG� ��ST��!>R|�FT���FT� FT� FPEMA�ILb �aA|p�FAULSHR�*��;pCOU_��q|pT���U�I< $d�S_�S#�ITճBUFkG�kG@�jpJ`p�0B�Tk�C�p�Rws�PSAV(e �R�+Bd�$ Cg�p��AP/d_ň�$̰_�Pec �iOT�����P@����jA�gAX��sq:p�P��\c_G:3
�YN_e!�pEJ0Df�W�r�d"UMO_0T��F�� �E2���^Јq	K��ey&^�5rH 8)�4��qL���nqL�S�cC_ܐ��K��pu�t��R�A�u�X�nqDSP�FnrPC�{IM5c�s�q�nq��U�w{0�0��PI�PR�nsN!D�@�sT!H��"ûr� Tߑ�s�HSDI�vABSC_�9@`�V��x�v���c~����NV��G ��~�*@�v�PF!�`ad�s0p�a��SC��\��sMER��nqF�BCMP��mpET��⌐M�BFU�0D�U�P?�M�B
�CD�yH��`�S9pR_N)O�ዑN� %�i�Xcg��PSf�C�@%v�C���a~Qd��`U OH����c  d�������}�锍� �9疗疢疮A*�7�8�9�0T��1��1
�1�U1$�11�1>�1K��1X�2f�2���2�
�2�2$�21�2�>�2K�2X�3f�3R�3��
�3�3$�U31�3>�3K�3X�94f��QEXT�TP <sK�p<6p��p2ǋ��QFDR^�QT�PV���b	2p�v�	2REMr�F��0BOVM�sz��A��TROV�ɳDT3`��MX��I�N��Q0�ʶIND����
	�i��`$DG�a{#��4P5�9D���RIV"�=2�0BGEAR�qIO�K��;N0p}ة��(���@�0<Z_MsCM@	1 �F|0;UR"�R ,t� a�? P0�?\��!?��EG ��`a��e�SG � 5P�a�RIM��@��SETUP2_ gT � �STD6� ��<����I�C�`��RwBACrU T[ �RTt)Nz%��+p�IFIQ!+p��А���PT{b[�LU�I1TV � Y�PUR�!�W2�r�<qv��P�� I��$��S��?x#�J�QpCOw`�cVRT|� x$SHO���SASSY��a?5P8�W����A�W�RKFU��15q��25q���*@�X |�N;AV�`��3����*@�R=1��VIS�IJД�SC���EP�c�\�AV��O���B%EX�$PO��I\ ��FMR2b�Y o�X�}p� bpNt�{ߍߟ߶ơP����_f�G�_���B��M4�Y�k�D�GCLFR%DGDMYLD��7�5!6H.�04%�MR�3SZ�@��	 T�FS�`2T[ P!��bs>�`$EX_��B�1�`Ā\2�3�M5��G��9\��
���PWeO�&D�EBUG��"��G�RR�spU�BKUv�O1�� 0PO� ;)' ��' �Mb�LOO�ci!S�M� E7b������� _E ] ��@Y� �TER�M�%^�%[�ORI�Bq� _�%1SM_OpL� `�%^���(�a�&�@UPRbg� -���]�#0^��G:0E�LTO{Q$US]E��NFIc1G2���!���$4_$U;FR��$j�A1�}0=�� OT�7��TqAX�p��3NSTCp�PATM�d@�2PTHJ�;�E4P_bD�H2ARTP`R5�PPa�{RG1REL�:�aS�HFT?�H1�1�8_�N�R�8��& � $�'H@a�q�B���b�SHI@�U�� JaAYLO��a�a����Y�1��~�J�ERVA�3H7�Cp�2�����E����RyC�~�ASYM.q�~�H1WJ[7��E ��1Y�>�U2TCp �a�5�Q=��5P��@���bFORCpMKT�z!:c��'"`&0�0w0�a� HOb�f�d Ԟ2��& X�O�CA1E!��$�OP����V�t �����P��P��`R�Ń�aOUx��3e���R�5Ie h�1��eo$PWRL�IM;e�BR_�S�4��� �36H1UD�_C�RBt]e7�$HSu!�`�ADDR2�H}!G �2�a�a�a��R��x�f H!�S����u��u
�u�SExv���!�HSH��:g $���P_�D�H Y�RrPRM�_��^HTTPu_i�Hx�h (*��OBJ���b��$�2�LE�3�s�i� � #�"�AB%_
�Tp#�rS�Px����KRL{iHITWCOUw�B6�L `�rQ��U�`��`�SS��JQUE?RY_FLAQ1�pQWR�N1x�jpgP&��PU����O���q��!t��/t����_�IOLNw�k(��� CJq$SL�L$INPUTM_Y$;`��P,���C̀SLA� l׀�(�$��C����B1IOgpF_�AShm}�$L ��w��8AِU� 4@�_1��݃��情@HY�1ǧ����a[�UOPen `l�ő2��� �������[`P�c;`��	������NqUJ�a�o � K�N!EaG4�v7F�Da��2�J7VpOQR$J8q�7�I_1z���7_LAB�1�P|����p�APHI���Q{���D�J7Jx�-��_KEY�� �K��LM�ONx�p�$X�R_���)�WATC�H_��C��D�EL�D��y����eq �@Р1V�@&�U�CT�R�3U�i��*l��LG��r� !#�LG�Z�Rࢵ�c��c���FD��I ����\!����� ���� e�Dqf�ce�c�e�ΰ�e�� e���@0J_@�ѐ1j��qʦ�F�A�xǒĞ�Cd(��SB����c��c���ΰ��I�����ƍ ̷ƞ�RS��0  �(ʀLNe�<sѐ���)��6�"��UosD��PLM�C�7DAUi�EAwp���T�u�GH�R1o��BOOw�t� C���`IT\���� 8������SCR���㖇�DI��Sw0HRGX ���z�d(��o���w�W�o�X��z�JGM^�MNC�Hl�n�FN�a�Kn��PRG��UF���B��FWD��HL.��STP��V�� X��Г�RS�HzP��w�CdD��1Rz�: :�^�Unq��9���H�k�����Gw�@( w�`������s�}�OC/ v��EXv�TUI��	I��7�C�O������<@���	$���<@��NOANqAo�A2� VAI����tCLUDCS�_HI$�!s�O��
�SI��S��IGN���ɳ��h�Tc�DEV�<�LL�A��_SBUI �uP�j@mT��$��EMr����]���*"	1vP�@j@ހ��~p����1�2�3�>��� 
0w �C��x�Q@5������IDXa$9 [�����֥1�STƐR��Y� <@   v$E.&C.+�pmp�=&P&����	1x L ����`��4@r�`Na��eENwp�dp��_ y ap7�}px	b���# �MC7��z �C�CLD�PƐUTRQLI��TT�94FLG )"0�Q53�DD�57�t�LD55455ORGT�8�H2_ȲF�8!s�D/r�#�S{ �� 	59�455S�PT0��0y0�4}�6RCLMCD@�?�?Iƀ�1pM�p�^���|�$DE�BUGGugQDAT�AY��T �UF�E��T)!��MI�6p�T} d@��R�Q��0DSTB��`� �F��HA�XR��G�LEXC#ES$R>��BMZ`��~� �B4���BSq*�����F_z@�H��S[�O�H�MJ;PTH�� &Pv��m��QMIR� �s � []R�WRCT��N}��VUO�ZA�ZL�RC�PQC��Q�`D��O��^�CURPX_THqG�P�`R`|1�o)`/d55R^`�`S<�P �B_FR@^�a\fZ_��^ddpG���* �!KH�� \���r�Fv$MBu�L�I�q�cREQUI[REG�MO�lO�k�fB�$ML� MG�� ap���`|��cB��ANDU�Sz��>�5�Z�9sD��Q�IqN�p��Q�RSMf�(Sx� �Q�!E]�q�RA'qPST� 7� 4�LO�P��RI ��EX�vA�NG��AQODA5QG���@$�QG��MFh������"���%&�2ТfSUP��%4QF `RIGG>�� � ��0�#�1��Ӫ#Q��$$���% #n�א~�א��rP��8wAZw@ETI9�~��Q2�M\p9� tV�pMD�I��)��� �DA�H�pu���DIA���ANSAW,��w���D���)�!O7��0�Љ �QU��VB�70�B�L�p�_V@�ъ ��C���sX@�b|�ٰ��P���v���Pƴ�KES�!���-$qB����� ND2FB���2_TX�$XGTRA�1����`LO�ЪЋ$RG��B�F�8Ҍ|�g�_���rRR2�E�0� #W�e�A�1 ?d$CALI�@2��G���2�RINܩ���<$R��SWq0"DᣫABC�x�D_J��a����_�J3�
�1SPHs�P��P�-�3,�(��?���\�J�l�4�2�1O8IM� �2CSKP":��~�Y���J���2Q��̵��8̵·�p_AZ�2h����ELg�FAOC�MP�s�1!I�RT�A)�Y�1�i�G���1�K�> Y�ZW�ScMG�܀�4JG� �SCLP�uSPH�_� �0����������RTERࠧ�ol�IN��ACz��|��� ��r��} _N�я������1j�4��?R� �DI��1�L�DHP3��ё�$V��Rs��>$v��p�1�������E�H ��$BEL�?w��__ACCEL��ؘ����P_Rـ� ҡQT!�*aEX2L6b��3���׀c@��.a�����36cRO
Q_�m�J�P�p�2�p`��_MG��$DDm�����$FW�0݀�Ӊ����~�DE��PPA�BN��RO��EE `���0±�YAOP���oa_��YPaPC��YY����1- �!YN�@A��7����7�M�A��ig�sOL�de�INCa���q����B�����AENCS��Á�B�Ѥ�,�D+`IN"I6b��<ހ��NTVEk���23_U�����/LOWL�#F�0��DF�D�`��ȯ ��`RC����MO�S� wT�PP�2��3P�ERCH  8OO`�� z�q�!��4!$��!�)b��A6b�L�tW����pF�
4TRK��!AY[�(cOQI��XM�p/�SQ�� MOMc��BOR�0���D��㣧d��⍠D�U��7bS_BCKLSH_C���@ YO`?����*N�>ĵCLALM���18�?P6%CHK0� >�GLRTY�������Ѕ|1܁_�N_UMzC�&CzC{��ܡ#��LMT)�_L �0ú$+��'E�-�  �+� ���%��>��C�L!4�PC��HI��`q�%C@8�{��CN_��N"C�6��SF�ѯ	V!�p!����U1��5Y8CAT�.SH�����?a����X�7aX�L�n�P�A�$��_P�%s_ ����Pn ��`rDc%aJAaPfC	 OGs7>�TORQU�A� Li���bd����B_W�IU�n��D_Ө�Ee��EI�KI[Ie�F�P�As�JX��w��VC��0�jS1�q^o��_��wVJRK�q\�R�VDB��Mt��MPp_DL_��GRV�D�T_��Te��QH_^��S�#j�COS0k1�0hLN �PSktUZd_�Uiv�Ui 'Q�jlEQ�UZN`d�QMY\a�h<b��Dk��iTHET0$N�K23e�rY�]`C�BvCBY�C��ASrqDr'TRq_�Rqv�SB_�pr*uGTSֱ��C0��qO�;C_�<�z�c$DU` ���r����xR�v���Q���53�NE��7�I�^`q#;��$=�qA�u;�D�"e-h-aLP!H0e����StU�� e���e��f�����f�=�V]�VR�O�u�V���V��V��V��V*��VɋV׉H]����|�t��1����H��H���H��HɋH׉OJN�O]�O�s�O��UO��O��O��O��OɋO�fF�?q���e��P�SPBAL�ANCEc�=1LE6�pH_uSP��pf��f�fPFUL�C������e��1=�+�UTO_[ �E�T1T2_���2N B!�������� ��p(�ҚӞT
O���>�@INSEG��=�REV��= ��DI�F3�1��1�1�&OB�&!�S��2�@��M!�TLCHgWAR��T�ABBA~�$MECHHq��`V�\�q&AXVP�4u�4�@�T�� 
pv��Ab���ROBn �CR���j2 ���MSK_֠�ԓ� P j�_�R ���2����51�2���������$��>�IN�ű�MTCOM�_C\P�Д  �h���$NO�RE��Q��.�@�7� 4�@GR�Ba��FLAű$XY�Z_DAQ����DEBU��f�.�m�� �$/�COD�! �҇b���$BUFIN�DX��B_��M{OR��� H�� ���E&��~�^�$޲���o1�� T=A������Ѱ�G�Ҙ � $SIMULp@�С�x�\��OBJE��>\�ADJUSz�m�OAY_I�A�D��OUT�@�Ԡ_�_[FIb�=��T�@ ��������q����������D,�FRI4��T�RO�@���E�A�OPWOܷP���,��SY�SBU+���$SO!PT���;!_�U^���PRUN0҅�PAB��D��`�Y� _��2z��AB��
0��/IMAG!����PϱIM���IN��P����RGOVR!D�v�e��P����� ��L_R�zA(�"��0RB� � 1MOC_ED��b� 
0�N+�MW	1�MY�191  �S�L����� ���OwVSL��SDI5�DEX�3��3
�	V�@�N��A��� ����n�C�0T���d�_SE9T�@��� @�@!��RI^���7_Lq@YL���x�.�0 ���Ta��@�ATUS�$T�RC���ҔBTIM��I��l41�sU ��� D��E���4�E���8� & �EXE�r! L� "�)�0��ƗUP��!IS��XNN��1ldQ^�	�PG>՟L�$SUB��V��ZJMPWAI2�0P��%LO� ���̰[�$RCVFAIL_C�i�!R��i�r�e1�0�4����%�`R_PLZD�BTB�A�2i�BW�D�&Y�UM�@�$I�G�������0TNL�0�$@2R'�T�~@�@<��PPEED5 �3HADOW�@c�Y��f�E��4�p!DE�FSP�� � L��|��0_�0���3�UNI����0C!R� L�`̰P�&p�P1�����Ю@@^Ѻ�� ���X�N�GKETB�@��	@�P42��� h �pSIZE�����ഒ�`ASx�ORZF�ORMATK�*4C�O~ \AǲEMn��|D�3UXC���PLI%2��� $�I�OMP_SWI�/��E��Wi�Js�!�P
0%0AL_ C��@�0"�gPBJ�DpC�D��$E�!�J3D�H�{ TV@PDCKC |m�X�CO_J3r��RQRĢ�	_] ���@C_/1A  �; �h�PAY�qҖ�T_1�Z2�S�@J�3�p�[�U�V�S6�TWIA4�Y5�Y6�MOM�c$cc$c4c;�B� ADcHf�cHfcPUSpNR )duecueb�2�A����` I$PI ��Ulq�U*s�Uus�U js�UUt�f�kit�t��v��v_!��m���:v3HIG�Cv3�% �4iv�4�%� ��iv�s�xx�!�y�!�%SAM�����tiw�s�%MO	V��$�'�
�ް)p %��� #��0�P2��P�%�0�5�`!��@��H��#�INj��@�sq� ��h��"s�������Ӌ�GAMMǦ����$GET���Є�D��T/�
z�LIBRt9!W2I��$HI8 !_��%�H�E"�U�1AO�r�c�LWJ��� ��r���c��Rn�M0�A�C50� a ?^I_�p2�/��B �X�AY��$c/�Hf���C �$,X W1���IXRk��D�>�A!�$@�LE@ �8q`���Xq��Z0_MSWFL�$M�@SCRI(7���)q��T"E@�A����P��UR�$�v�K�S_SAVE_DX-B�;#NO�PC` <"�TB�&��_�a�YW� �i�Y�`����pkR#uܸ�SD��p#�s0� @�,�$�cxY�svY�x�@�<����<!!�@M��ũ � "�YQL�c��Y��S�� 6�0�� 0����J��� �����	�t�Wq���A�`��1�t�M����CL���Q��o ��1T"�@M3�*� ό $��G$WRГ����QR�oT P�vTP�}TP�T0���+��C;�@X�0O�~S�AZ�տ@��Uԫ[ �ՑOMK��V���������̿`CO�N�� �c�Q_v"� |=Q�B�$i��c ��cB��Z���j�A� ������t�P��P_A�PM� �QU�p � 8�@QCOUM�i�Q�TH/0HO��G�H�YS�@ES�F�U�E2�8�E@O�D� � �@P0�@�`UN����q�OVr�а P����%$��W2�ROGRA���22�O����IT�����t�INFOXѱ ��A�����p�O�I� ((�SLEQZv/Nu/ �����OS��s$� 4�@ENAB~�� PTIONZ�4(r�\�4cGCFl�0�J� �A���,�R�����OS_sED� �е �NR��K�:G�E��sNUAUT^�COPY�8 7�1j�MN�NAEPRUTf� HNֲ OU�B�0RG�ADJXѶTBX_t��2$�0��мW�P����v3���#EX� YC~�^DARGNSh����ޠLGO��PNY�Q_FREQ�bW`��MvM!�D��LA���D!�c��@CRE�3�R���IF�a��NmA�q%�$_G}4�TATB0�$>�MAIL�r2��!��B��1x�!1�$ELEMl� �s0vFEASIy@���@��2@@K�66�V�2�I���0�D"8qJ��k2AIB�APE��vpV�!�6BAS&R�52��aqU�p��W�$�1~�7RMS_TRe3 �A���3�ӓp�r�!�4c + !"������	B2 2�  ���ԇ�(F�2'G�2/��_����2SG�g��DO�U��N�!"PR�e�m �6GRID���b�BARSZwT9Yz�"OTO?`X�W� ��_�$!���B�DO��i� �s ����POR���C�f�BSRV� ),TVDI`�T�P0Q�CT� MWCpMW4KY5*KY6KY7KY8/Q��F�l��$VALU�35�(4��}Fh�� u�Y����C�!2�� AN4��R�!RR!2�TOTAL�s�a2c�PW:#I�AHdREGGENFj[b��X�8`��R%��V-�TR�3�rFa_S8��g[`�AV���b��2E�#��@L�1�-cV_�H�@DA-��`pS�_Yf���^&S�A�R-�2� �IG_SEC�`R�%_���dC_�F�Q�E��q�OG6�kjxSL)GEpl�� >�_%���/�0`9`S���$D�E.QU>����sTE|���P�� !�a���aJ�v^�3IL�_Mm$;����`��T�Q-�6���0Ƨ��V�h�Cv�P�#1��M���V1��V1��2���2��3��3��4��4��$��`ӓ%�� �0����INA�VIAB=�p�]��d�2`�U2l�3`�3l�4`�4l�X�WB �pB�����D $MC�_FP���%�LPC�B�f#cMo�I��oC ��6��q���KEEP_HNADD�!#��0-�	C�ѫ C��A⒤�D�O&�"�{��3�D���!a#D�REM[�@C�8a�B������U�$�eC�HPWD  �#�SBMSK~�BCOLLAB/���P@�$a�" IT�$ ��fȕ��� ,�(�FL{�W�M�YNTڐ1�M��C`r�G`�UP_DLYX���DELAc�9a�"�Y�AD-��AQ�SKIPw�� �4P��O��NT9�����P_������ ��÷�aѹ�ѹdPк qPк~Pк�Pк�Pк��Pк9��J2RT ���qX�0TG# r���qr�� �r������RDCS�� �_�R�R1�o�=��R�!��J��*DRG�E� T3�ÆBFLGp'����*DSPC���!UM_r�!�2T�H2NrA<�e� 1�  ��@v� 11��� l��0��O�v�ATy�� .��Q&�������� �*D�Ҙ���H��� +_U�2]��c�u�p�ߙ߽߫� U�3]��������(�:� �U�4]�� ]�o�����V�5]���������"��4� U�6]�� W�i�{������� U�7]��������
.F�8]��Qcu������S�L�R��1V�p`�L㙠-E%$рp�eL)fcIO��I��R��POWEC��� M0��� �T�#d �+��$DSB] � �""c^�QCB��R��M
E�+�R�	D��0E�"���MD"'��M�E� yD�p�'DBG_~@aPD�3%!eaPG
A�@���@S23�2i� ����<P��pICEU�2!`<k$�pARITq!a�OPB�rFLOW>pTR(.b��@�qCU� M%3UX�TA�qINTEORFAC�$��U`���SCHA׃ t�ݐ"!hp��$�`�`OM'p�sAD���0Iᓴ0Q@A+��TDSv`���8c3�EFA����r�S� k��`8b� q��R H��6A �ٶ�q  2�� �S��M �	O� �$)�s�0��
eC2`_%pFDSP)FJOG�`�#�p3_P���"ONg�u���'�	6Ky0_MI1REAb$wpMTY��CAPK�wp4Ц@�4"A�Sp}@r"At �EBRKH<16=��R��! �B�s�BBPo0�b<C@BSOCF��uNUD1pY16���$SVi�DE_�OPGtFSPD_�OVR�k��DLTRWCORbW� N�PbcVF�@�WB@OVEECSF�Z^p�S,rF�V� t'�UFRA�ZTO�$LCHa�u�2�#OVST��B@WQ����BCZ� r&PQ@]s ; @�TIN�``!_$OFSC`C�0@�WD|QdxQ%Q�,�E?PTR�!e"�A�FD���AMB_C��bB5@B<��!q�b�a�cSV��L�k0ȉ�s��RG�g�HAM�tB_=0�e-b_�M�`2�:`T$SCA8@�D�B?p�HBKo1~6TqIO��cu�pqPPA Wz�qhy�t{uu�:bDVC_W R#�p1 ��p���Q�u���x-s�u3�v3`��{�0p@�SQUR#7@~CAB ���,Ӟ`���`�h9��O�`UX~6SUB'CPU�O@S��� ���dp0ݱ���c�d�~��$HW_C]� �0ݱrpʆ�� �NÐ�$U��D��>�ATTRI�0���O@CYCLw�NE�CA)��CFLTR_2_FI�/����LP[KCHK�ՠ_SCT�CF_��F_�|��FS8��b�CHA��d�p���b�"��RSDU�`�Q�3��_T�h0Y���c� EM"��EM�CT��ݰĀ�����2�DIAG5R�AILAC�sx�M���LO	P7�/V����3� H�3��sPR��pS+� 90��C��q� 	,cFUNC:��1RIN���a$D����!ʰS_"@*?p䣸�Mt����MtCBLȰ���A0�
��
�DA�@�O���LD`0GPpq�w�*A�|�w�TI�����AĀ$CE�_RIA��AF�Pn#ò%`ȵT2bd�C}3�r�aOI��fDF_LY�Rl1��0LM`#FA  H�RDYO�AM`RG�|�Hސ�Q� W��MULSE��3��8P.�$J_ZJzR�W��[FAN_ALMsLV�#��WRN��HARD�@o6���2$SHADOW  `������V���!�Q��E_`s�AU��R���2TO_SBR ��6@(�逺sá@�_MPINF8`��8S�m�^�REG���DGy�K�Vm0��F�DAL_N�dFLۅ9�$Mm�l�D�hg O`L�K$g$Y("V1	�2~#�� ��CCEG[CGP
�A �~/U28S�;��EA�XE,GROB)JR�ED)FWR  �A_i�SSY�@D��@��S��WRI  �ɀ�ST�*C0�@nPE��&�w� �"@B���9a��5k�pOT�On�%`ARY�)C�e��,[@FI��@pC$LINK��GTH2��0T)_��9a%�69R[�XYZo2e�7s�OFFA`2� \�N�uOB'@����a� h0��FI���0�4?T��AD_J�!�2@lR?�pq������89R � ��	T�AC��F�DUWb$�9x�TU�R��X��z!�N�X��� )FL[��PH�0�� |���309ROa� 1�KN@Ms�/U3��{�������W3ORQ�6A��(��{��@O��N��Hp�34A��]OVEd("M00J��~��~ ��}F1|J�|�{AN��5�~ȱ)!e }@���ve�%0��%�6AERSA	|�E �`��E$A�Ā��ܥ��V�S�V�AXc�2V�� ҁ4�%8��)b��)w� �*�*r�*��*: �*q �*1� �&��) ��)��)��)��) ��)�9�9�'9�D189DEBU���$����0��1VbV�A!BV�Tq|Q^VIp�� 
B�s��+E�� 7G8Q7Gw�7G�7Gr� 7G��7G:7GqδF �Ȳ4��LAB��8)���sGROB�)��2pB_�,&�� uS��%��FQ*U�VAND� |�:$3�_�=!�YW 2qZ�^�`mX�|X5�^�NT��
c�PVEL���Q�T��V�SERVE��P��� $���A6�Q!�PPOHb����`��QN�R�����  $bT�RQK�
 ct�
`ߌgȲ2�e��Q�_ � l���a��'ERR��m"I� �P��raTOQ��L�H�$��f�G�U%�H�f��T��X� � ,�Q#e=`��R�A�a 2� d��b{s��d` ���$r����"��dOCG�p� � dkCOUN�T�� ��SFZ�N_CFG	a� 4ƀ��;�T�Ŀ����3�����b!qTq��� �(@M��o���`#������uFA���ö�sXd��{�y�aH��S��TO�d�PJ���PHEL��Yr�� 5k�B_B;ASf�RSR�֤�E^�S끐�M�1�g�M�2p�3p�4p�5*p�6p�7p�8�g@��ROO��`9�]�NL��LAB�SN�N��ACKFINpTo���$U��M��� ��_PUV���b�OU�P̠��-��f������&TPFWD_KcARwa��f`RE�T�,�P/�]��QUE����eU �����I ��C-�[�[��Py�[�SEM3A�AAH�An�qSTY�SOސ	�DI�ɠ}s���'���_TM��MANsRQL�[�ENDZ�$KEYSWI�TCH^�s�.�ĔH}EU BEATM��PE�LEvb��@J��Ur�F�s�S3��DO_HOMưOl���EFA PR��Prv����C��O8�<c`�aOV_M����IOCMG˗?�b.�HK��� �DX�׍pU�¹�M�����HFORC���WAR(�7P,�O}M� � @�4T���U��P3�1��2��3��4=��bp�O��L����b��U�NLO9����E�D��  QpNPXw_ASZr� 0����Ѝp��$SIZ���$VAP�eM_ULTIP��.��ŰA��� � �$H�/����B�S�}s�Cr`��FRI	Fm"pS��������{NFO�ODBU�� ~P�������U)�N��з� xU`SI�bTqE�8��SGL*�	TA� &opC��C���+�STMT�\�P���BWe,�SHsOWd�n �SV7 �_G�r� : $PaC�@p7#�!FB��-P��SPːA�����`VD�Оr�w� �WaA00^T ��ɰ��Ӱ��ݰ��簪��5��6��7��8*��9��A��B�ٴ� �׳A��y���F��70T���1�1"�1/�U1<�1I�1V�1c�U1p�1}�1��1��U1��1��1��2��U2�2�2"�2/�2<�2I�2V�9 ���p�2}�2��2��2
��2��2��� `�>`"�3/�3<�3�I�3V�3c�3p�3�}�3��3��3��3���3��4k	4�4��4"�4/�4<�4�I�4V�4c�4p�4�}�4��4��4��4���4��5k	5�5��5"�5/�5<�5�I�5V�5c�5p�5�}�5��5��5��5���5��6k	6�6��6"�6/�6<�6�I�6V�6c�6p�6�}�6��6��6��6���6��7k	7�7��7"�7/�7<�7�I�7V�7c�7p�7�}�7��7��7��7���7��p��P��Ub� `{@e��
�PV���Q�U��PR��CM�p�bMb�PR9` ��TQ_+p�R�P�e(a~��SQpY�SL�`�P� � L��jw��A�ؠ; xѠ�D��VALUju�%�x��A6XF�AID�_L��^UHIYZI~��$FILE_L���Ti�$��`�CS�Aq� h ��pVE_BLCK��RE��XD_CPU�YM��YA�us�_�T�w@Y*�F�R �? � PW-p�l�<aLAj�Sq�AcRaKdRUN_FLGde@dhaKdv�ke�a@d�aKeHF�Wd�`�Kd$PP�TBC}2�u� � �Bk`(���pĠ���dN	�TDCk`|r�b0�p��
u�gTH	�%s�D1vR��ESE�RVE��Rt	�Rt3���`�'p ��X -$}qLEN`���t	�}p)�RA����sLOW_�Ac14}qvT2�wMO�Q�	S���I.��B�Q�y��D}p�DE���LgACE,��CCC��B��_MA2��J� �J�TCVQ�r� �TX�s����������H�� ���J+���Mۄ"~�Jw������ ��q2�������6�JK(�VK��:�0>�:�sq/�J0O�>��JJF�JJN�AAAL>�t�F�t�n�4o�5/sX�N1����d��N��DL�p_XѩQ���aCF6�� `�PGROUDPF�Q����N�`C�� �RE�QUIR=rؠEBqU��yq܆$T��2�6�zp ��$$�CLAF� ���ݐ��*�*� qO���X�e����k�IRTU�ALW�i�AAVM_WRK 2 ��� ?0  �5a�ͯr٨ʯ�� ��A	s@�3�*����!�^�E�c�������`��ɿۿ㴧�BS�@��� 1x�� <��(�:�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�� �����������
�� .�@�R�d�v������� ��������*<8�~pN�LMTu�?���  dQI�NZlPPRE_EXE}� �~A�AT�ʖ���IOgCNVՒ~ �h�P�US���I�O_�  1��P $���I�4��1��?�?_ Tfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(��:�Q LARMRE?COV �c��LMDG �(BLM_IF m? ������+���N�`��r߄ߕ�, 
 �߾�9�E��������ANGTOL�  �
 	 �A   Y�k�Q P�PLICATIO�N ?�� ����ArcT�ool �� 
�V9.00P/0�3j�+�
883340����F0����1612�������7DC3��+���None+�F{RA+� 6��LP_ACTIV��	j��UT/OMOD� �Ո	�P_CHGAPO�NL�� ��OUPLED 1�  !3���CUREQ 1�  T=	=�=	�������=_ARC� Wel=�A�W�ՕAWTO;PK�HKY�D y�9'EK ]o������ 5/�/#/A/G/Y/k/ }/�/�/�/�/�/1?�/ ??=?C?U?g?y?�? �?�?�?�?-O�?	OO 9O?OQOcOuO�O�O�O �O�O)_�O__5_;_ M___q_�_�_�_�_�_ %o�_oo1o7oIo[o moo�o�o�o�o!�o �o-3EWi{ �������� )�/�A�S�e�w����� ���������%�+� =�O�a�s��������� �ߟ��!�'�9�K�`]�o����OTOC������DO_CLE�AN�����NM  H���^�p��������A_DSPDgRYR���HI��<�@M��&�8�J�\� nπϒϤ϶���������MAX��������
�X�������PLUGG�����
�PRC˰B:�"H����d�Oi�Կ��SEGF��� �� ����:�L��&�8�J�8\����LAP�� ��������������"�4�F�X�j�|�q�T�OTAL,�U�USWENU���� ߨ����O RGDIS�PMMC� ��C���@@M��O���߹RG_S�TRING 1~��
�M���S��
__ITwEM1i  n�� ������� '9K]o������I/�O SIGNAL�cTryou�t modej�Inp Simu�latednO�ut-,OVE�RR� = 10�0mIn cy�cl!%nPro?g Abor7#n�$status��${ cess F�ault�,Ale�r�$	Heart�bea�#�Hand Broke� ��/??%?7?I?[?m??��e��w �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O��O�O__�?WOR ��eKQ�?%_s_�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�o�nPOc�!�`c[ �o$6HZl~ ��������� �2�D�V�h��bDEV�n������̏ޏ ����&�8�J�\�n� ��������ȟڟ���>�PALT�=7� c_�_�q��������� ˯ݯ���%�7�I��[�m������%�GRI�e۱O����� '�9�K�]�oρϓϥ� �����������#�5�G�ɿ��R�=��Y� �߹���������%� 7�I�[�m������������m�PREG ;�$����K�]�o��� �������������� #5GYk}����$ARG_KPD ?	������  �	$�	[��]���� S�BN_CONFIQG� �%!$"�CII_SAVE  �D;� �TCELLSET�UP 
�
%  OME_IO���%MOV_H8���REP�����UTOBACK�s�	AFRwA:\� �,�^'`� �<(�� M+@ �23/04/�01 14:33:48���/0�/�/�/-,��?/?@A?S?e?w?�?��? �?�?�?�?�?O�?5O GOYOkO}O�O�O,O�O �O�O�O__�OC_U_�g_y_�_�_�_�Ё � (!_#_\AT�BCKCTL.T�MP DATE.D:��_oo,o>o#�INI:�o%7~#MESSAGS�]a^� hkODE_AD�V7G�eO����o#PAUS�a!��� ,,		�� ��ow �o-9;M�q ���������;����d�`TSK�  �m</Bo UgPDT�`[gd����fXWZD_ENqB[d3��STAZe�����WEPLS�CH R+   b��.�@� R�d�v���������П �����*�<�N�`� r���������̯ޯ�����RODނ2.�4���/��>� %V�{������� ÿտ�����/�A��SϾWEROBGRP`��r�GWEWEL �2�D� ��h�����'�9�K� ]�o߁ߓߥ߷��߼	�XIS%UN��8�D��� 	r�� ��@�+�d�O��s���������MET�ER 2b�_ �P��&���J���SC�RDCFG 1v�! �[[?�������������5/�
QW��M_ q����2� %7I���!GR�Р��o��PNAME 	��s	$�_EDY`�1s�� 
 ��%-�PEDT- v��/*/j�������.��µ���X��/:����%2�/ ���/a/��G(�//?v/�/?�/�#3g?�/�? �/>�?�?B?T?�?x?�#43O�?�O�?>\O@�OO O�ODO�#5�O oOL_�O>(_�_�O�O�__�#6�_;_o__ >�__o�_�_No�_�#7�oo�o+o>�o+ ro�o�o�#8c/�//�=��>P�t�#9/��|���=X�Ï
����@��!CR�/�oG�Y�} "���ԏ�|�
���?NO_DEL���GE_UNUSE���IGALLO�W 1��  � (*SYS�TEM*��	$S�ERV_u�.�G�P�OSREGP�$8r�.�G�NUMu������PMU����LAY��.��PMPALTǧCOYC10Ԟ�Ѡ<ծ�ULSUǯ����r���L#�\�B�OXORIy�CU�R_I���PMC�NVæI�10�����T4DLIB�@�b�	*PROG�RAO�PG_cMIծ���ALߵ����B<�G��$FLUI_RECSU�u��j�������������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r�������������e��LAL_OUT 6��q#�WD_ABO�R��i�ITR_�RTN  �����l�NONSTO���� ��CCG�_CONFIG �7�7���8������E_RIA_�I���, ����FCFG ����5_LImM^�2� � 	n���<�j�ߥ蜀�dP}AV�GP 1?��-�?�C�� C��  C�b�fԪb�f�f�b��f0�D`�DD���
��4���Dv�DZlT~����Vx�D/�9�C��M�W�a��?����HE��u�"G�_P��1�  ��d/v/�/�/�/��/�/HKPAU�Sf�16�,  ���/ ?6�?L?2?\? �?h?�?�?�?�?�?�?�O�?6OHO.OlO
O�9?��h�CO�LLECT_90s	`�N�GEN߰���~��B�ANDE�C�s���12�34567890�!W��a�O_1V��
 H+���)l_�_a� k_}_�_b��_�_o�_ �_	obo-o?oQo�ouo �o�o�o�o�o�o: )�M_q��@�����Fm�K� �N�FIO !
Y�A��������ظ�ʏb�TR� 2"F�(��}�
�؎���#q�� %[�_MkORm$� �) ���������ǟ���Pٛd��n%r�, %I?	!	!�>���KH�*��$R9&�Ow��v�v�C4  A�l�
� x��AA��Cz  B�fPB}���C  @��������:d�U
\�IS'f�\��T_DEF*� ��%�+�����IN�US�&,@�KEY_TBL  ��,v� �	
��� !"#�$%&'()*+�,-./*W:;<=>?@ABC��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~�����������������������������������������������������������������������������������������������������������������������������������������6�d�L�CKI���d�I�ST�As�>�_AUTO�_DO��m���I�ND�D�δAR_T1�Ͽ�T2��������A�XC� 2(�q�cP8
SONY XC-56{��u��U��@����� ��А~�HR5XY ���έ�R57����ACff���6�H� $� m��Z�������� ���!���E�W�2�{�܍��TRL�LE�TE!��T_S�CREEN ~�
kcsc"�UD�MMENU �1)�	  <u��1�:o `CLr����� �� &_6H �l~����/ ��I/ /2//V/h/ �/�/�/�/�/�/�/3? 
??B?{?R?d?�?�? �?�?�?�?�?/OOO eO<ONO�OrO�O�O�O �O�O_�O_O_&_8_ ^_�_n_�_�_�_�_o �_�_oKo"o4o�oXo jo�o�o�o�o�o�o�o�5+���_MANU3ALH��DB9�0������DBG_ER�RL�*����C >���~uq�NUMLIM���dn�ޠDBPXWORK 1+���L�^�p�������DBTB_�� Q,�}����u�RqDB_AWAY}s�͡GCP n�=s����_AL
����yrYGл�n�nx�_�p 1-q�
́.�
;�y�z�g�l����_M��IS�����@A���ONTImM���n��ޖ�4�
X�I�MOTN�ENDM�H�REC�ORD 13��� �����G�O� t�b���������į֯ m�ޯ�t�)���M�_� q������˿:�� ��%���Iϸ�m�ܿ �ϣϵ���6���Z�� ~�3�E�W�i��ύ��� �� ��������z�/� ��:���w����� ��@���d��+�=�O����s�^�l�����Oi������b�M��sN��������[���);�_JX���W�����N/��9/�k0�.:/q/�/���TO�LERENC��B��>��L��upC�SS_CNSTC�Y 24,���p�/<���/??(?>? L?^?p?�?�?�?�?�? �?�? OO$O6OHO�$�DEVICE 25�+ І�O�O �O�O�O�O__+_=_�O_���#HNDGDg 6�+ՀCzi^_LS 27�Ma_ �_�_�_oo'o9oc_��"PARAM �8U�%�duKd�$SLAVE 9�]�nW_CFG :�koKcdMC:�\� L%04d.'CSVJo<�c�ofr6+"A sCHp�QA��Kn*_}g�Kf�Or|q�zyyq�`�JPѬsk~<�ρ��lRC_OUT �;�MρOo_SG�N <K�4����mE08-A�PR-23 11G:15p�a/�13��4:3?��F V�t�g�c�Knd��+�@�S�Þ��j�x�z��cV�ERSION ��V4.0�.1��EFLOG�IC 1=�+ 	�x�`��q���PROG_ENqB)��V2�ULS�� �V�_ACC�LIM����c�q�WRSTJ�Nɐ�3��a�MO�;�uq�b��INIT� >�*K��a OPT�` ?	��Ȓ
 	Rg575Kc�74!�56"�7"�50F�ׄ�L�2"��xp�އ��TO  �z�ů߆]V֐DEX��d&���pݣPATH ;A�A\˯*��<��+HCP_CL?NTID ?�c �{G#|��!�IAG_GRP {2C�i Q�	��ؿÿ��� ���Dϒ�mp1m�10 8901234567n���=�� ?ϜϮω������r������!� 3���\�n����q� Gߩ߻ߙ�����{�� ��9�K�)�o���U� g������������� 3�Y�7�i����+�u� ��������/ gyW��9�� �	�-?�>� �:ϫ����|�@��;/&/_/�˰_O 4Q/�/A/#�/g �/?!?혒$-?W?�/ g?�?o?�?�?m�?E/ O�?ODO/OhOSO�O wO�O�O�O�O�O
_�Op.__R_��<�p c_�_�_C_�_�_ �_�_�_o0o�_@ofo�Qo�ouo�o�o�o��C�T_CONFIG� D��ʓ]��eg�u��ST�BF_TTS��
@J�)s��}�xq<v�p�MAU��?�Q�MS�W_CF�`E�� � ��OCVIE�WPpF�}�a�� ������*�<��� �e�w���������N� �����+�=�̏a� s���������͟\�� ��'�9�K�ڟo��� ������ɯX����� #�5�G�Y��}����� ��ſ׿f�����1�XC�Uϡ|RC�sG]r!�c΍��ϱ������
���.�tSBL�_FAULT �H�ʥxH�GPMS�K2w[��`TDIAOG Iy�qUt���UD1: �67890123C45��x��c�P�o ����*�<�N�`�r� ������������(�;�Vp���@8r��|\��fTRECP����
�ԣ��������� ��1CUgy �������	�0�B�?f�UMP_?OPTION2pT�FaTR�r3sX���PME1uuY_T�EMP  Èϓ3B�Vp��A��UNInp4u����YN_BRK �J��bEDIT�_y�ENT 1K~��  ,&�`R/P@/}/P�l/ �/�/�/�/�/?�/'? ?K?]?D?�?h?�?�? �?�?�?�?�?�?5OO YO@OhO�OvO�O�O�O �O�O_�O1_C_*_g_�N_�_r_ MGDI_STA��q�%�NC�S1L�{ ���_�_P
Pd 7Yoko}o�o�o�o�o �o�o�o1CU gy������ ��� �.�Fa.�T� f�x���������ҏ� ����,�>�P�b�t� ��������6����� �#�=�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��۟���	��5�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹�ӿ���� ��-�#�I�[�m�� ������������� !�3�E�W�i�{����� ������������7� ASew���� ���+=O as�������� �///9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? �?�?��?�?�?O'/ 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�_�_�_�?�_ �_�_oOo;oMo_o qo�o�o�o�o�o�o�o %7I[m ���_����o )o3�E�W�i�{����� ��ÏՏ�����/� A�S�e�w������� џ����!�+�=�O� a�s���������ͯ߯ ���'�9�K�]�o� �������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߷� ����������-�?� Q�c�u������� ������)�;�M�_� q������ߝ������� 	���%7I[m ������� !3EWi{��� ������/// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?���?�?�? �?/O'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �?�_�_�_�_Ooo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu��_��� ��_��)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� �����ǟٟ��� !�3�E�W�i�{����� ��ïկ�����/� A�S�e�w��������� ѿ�����+�=�O� a�sυϗϩϻ����� ����'�9�K�]�o� 鿛��߷��������� �#�5�G�Y�k�}�� ������������� 1�C�U�g�y��ߝ��� ��������	-? Qcu����� ��);M_ q��y������ //%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?i?���? �?�?y?��?OO/O AOSOeOwO�O�O�O�O �O�O�O__+_=_O_ a_{?�?�_�_�_�_�? �_oo'o9oKo]ooo �o�o�o�o�o�o�o�o #5GYk�_� ����_���� 1�C�U�g�y������� ��ӏ���	��-�?� Q�c�}��������� ɟ���)�;�M�_� q���������˯ݯ� ��%�7�I�[�u�g� ������ϟ����� !�3�E�W�i�{ύϟ� ������������/� A�S�m���ߛ߭߿� ٿ������+�=�O� a�s��������� ����'�9�K���w� ���������������� #5GYk}� ������ 1CUo�y��� �����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?g U?�?�?�?��?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_�!_3_E__? �$E�NETMODE �1M�5��  o0o0�j5�_�[nPRROR�_PROG %�{Z%i6�_�Y�UTA�BLE  {[��?-o?oQo_g�RSE�V_NUM �R?  ��Q�`��Q_AUTO_ENB  �U�S�Tw_NO�a N{[��Q�b  *�*�`��`��`��`�`�+�`�o�dHI�S}cm1�P�k_AL�M 1O{[ �2j4�li0+�@�����_vb.�`  {[�a�R�2�nPTCP_VE/R !{Z!�_��$EXTLOG_7REQ3v�i���SIZ���STKڪ��e�TOoL  m1Dz;r��A �_BW�D�瀠f��R��D�I� P�5���Tm1�STE�P)�;�nPU�OP_�DȌlQFDR_?GRP 1Q{Y�a�d 	-�ʟ�P����E%�ڭ�?�#��[���� �
� ��������!�� D�/�h�S���w���������ѯ
���.��W
 $�]�fvM��������ޫ�B�  �A�?  @�33��UO��Ϳ��9��$�F�6 F@�]�[�g�"σ�F� �?�  �Ϙ�<P����;O��9� n���r���r���i"I��������:��q!�s�[FE�ATURE R��5��QArcTool D��m2Engli�sh Dicti�onaryO�4D� Standar�dH�Analog� I/OG�AZ�e� Shift��r�c EQ Pro�gram Sel�ect��Soft�par����Wel�d��cedureys��@�Core���?�Rampingn��uto��wa'�UpdateM�m�atic Bac�kupM�{�gro�und Edit�E�R�Cameraz��F��Cell�����nrRndIm����ommon �calib UI�����sh�����c�&�.���neC�.�t%y��s����n���Monitorb��ntr>�eliayb��N�DHCPD����ata Acq�uis���iag�nosw����oc�ument Vigewe���ua#��heck Saf�ety	�R�han�� Rob��rvB��qF
�N�ks" �F��(�R�xt w�eavx�chJ�x�t. DIO$�nsfiG� endS Err��L��%s�	r���  �L��FCTN Men�u; �  TP I�nfac(�R�G�en��l�Eq �L�]��p Ma�sk ExcO g�HTJ��xy �Sv#�igh-wSpeS Ski������$�mmuni�cv�on�Hou�r1����Mco�nn}�2(ncr�Lstruc�M�K�AREL Cmd7. L�ua�E#�Run-Ti� E�nv;(_�+z�s�x�S/WO�Lic�ense5"� B�ook(Syst�em)L�MACR�Os,�/Off;se�MMR�����MechStoEp��t�����%i����6xS ��x�1>od��wit�T8�����.$�r;Optm8�?�#��fil"�'�g��%ulti-�T�E�P�PCM 'fun4'�9o��6�E�MRegi� r,��6ri F
KRF���Nu����nH��Adju�hN�Ҵ٦MtatuNA�O
QշRDMUot`�s�covei��Eem0�nw��ERZ� N^ues��9Wo$��_0N�SNPX b�"H�SNJCli}^��urhӝ_z�Q %4ujUo� t1ssagE�jU�A��{_F� U��!n/I|KeMILIB;o~bP Firm^�:%nP1Acc�����TPTX��del�n� XoaA��%&mo�rIP SimulQa����fu� P]��j���3&��ev�.eV�ri3 �o?USB po����iP� a bunexceptS P(DXbu�uVC�r��8V���rvo�u�[��{S�PSC�e
�S�UIK�W� �8<�b Pl�FX�Z�� �M�#�FQ�xuvn�ԇGrid
Qplay΍"`��eR�r.wڊ�RC��g�100iD/1�450��larm Cause/P�edj�Ascii���Load" v�U3pl����yc��k"0Y@Pp@ %RAp��<l�"�NRTL�oS��Online Hel���6L�6L@IA��trG�64MB� DRAM��\�F�ROe���tl!�0.�L�mai#��[�L%�Supmr�1NIР� �cro�LS�U���V�Rmi܉�vrt2SK������W� i�������̿ÿտ� ���%�/�\�S�eϒ� �ϛ��Ͽ�������� !�+�X�O�aߎ߅ߗ� �߻���������'� T�K�]������� ���������#�P�G� Y���}����������� ����LCU� y������� H?Q~u� ������// D/;/M/z/q/�/�/�/ �/�/�/�/	??@?7? I?v?m??�?�?�?�? �?�?OO<O3OEOrO iO{O�O�O�O�O�O�O __8_/_A_n_e_w_ �_�_�_�_�_�_�_o 4o+o=ojoaoso�o�o �o�o�o�o�o0' 9f]o���� ����,�#�5�b� Y�k�������Ώŏ׏ ���(��1�^�U�g� ������ʟ��ӟ��� $��-�Z�Q�c����� ��Ư��ϯ�� �� )�V�M�_�������¿ ��˿����%�R� I�[ψ�ϑϾϵ��� ������!�N�E�W� ��{ߍߺ߱������� ���J�A�S��w� ����������� �F�=�O�|�s����� ��������B 9Kxo���� ���>5G tk}����� /�/:/1/C/p/g/ y/�/�/�/�/�/ ?�/ 	?6?-???l?c?u?�? �?�?�?�?�?�?O2O )O;OhO_OqO�O�O�O �O�O�O�O_._%_7_ d_[_m_�_�_�_�_�_ �_�_�_*o!o3o`oWo io�o�o�o�o�o�o�o �o&/\Se� �������"� �+�X�O�a������� �����ߏ���'� T�K�]����������� �۟���#�P�G� Y���}��������ׯ ����L�C�U��� y�������ܿӿ�� 	��H�?�Q�~�uχ� �ϫ���������� D�;�M�z�q߃ߝߧ� ������
���@�7� I�v�m�������� ������<�3�E�r� i�{����������� ��8/Anew ������� 4+=jas�� �����/0/'/ 9/f/]/o/�/�/�/�/ �/�/�/�/,?#?5?b? Y?k?�?�?�?�?�?�? �?�?(OO1O^OUOgO �O�O�O�O�O�O�O�O�$_Q  OH541S?Q2DVoR782EW50EUoJ614iW76EU�AWSPQW1�WRkCRuX8�VTU�V�J545iX�VVC{AMEUCLIO�V�RI�WUIFQV6��WCMSCh�VS�TYLiW2�VCN�REQV52�VR6�3PWSCHEUDO�CVqfCSUEUO{RS�VR869iW�0tW88DVEIO�fR54\VR69��VESET�W�WJ�YWMGEUMAS�KEUPRXY5h7&EVOC�V�`3�X\VX�`hXgX53�fH^xwLCHvOPLv�J50HvPS�wM�C�W�p�g55tVMgDSW�w;wOP;wMPR�Va`0v�`hVPCMg0��`tW�50�51�W51�P�0�VPRS�g6�90vFRD�VRMsCN)f�hH93hV�SNBAg_wSH�LB)fM߇a`XgNuNlx2hVHTC�V�TMI4fYP�fTP�AfTPTX�EL���p�g8[WYPDVwJ95�VTUT<w�950vUECvU�FR�VVCC��O�VVIP4fCSC�L��`I�xtVWEB��VHTT�W6WgW�IO��CG�IG��IPGS=�RC�4fHZXR66�VRU7�gRN�2HvRjz�40vu�tV`DVNV�D�fD0��F�C�TO�WNN0vOL�'hENDQVL×S;LM�fFVRe X K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩπ����������'��  H54�1)�C�2H�R78�2I�50I�J61�4y�76I�AWSuPY�1��RCR���8��TU��J54y5yܘ�VCAMI�oCLIO�RI��UIFY�6��CM�SCY��STYLzy�2��CNREYڻ52��R63X�S{CHI�DOCV��wCSUI�ORS�گR869y�0��8�8H�EIOh�R5�4h�R69��ES�ET�۷�J��WM�GI�MASKI�P�RXY��7I�OC(��3��hڅ�x�w��53�HLCH��OPL��J506��PSgMC��u ���55��MDSW���OP��MPR�(�����%�x�PCMbH�0����50[51��51X0�ڷPRSx�69��F{RD�RMCNy���H93x�SNByAI�SHLBy�M+���NN(2�x�HTC��TMI���e��TPAh�T7PTXi*EL�u ��8g�e�H�J95n��TUT��95��wUEC��UFR��VCC8<O��VI�P��CSC�*��I�i��WEB��HTuT��6��WIO�:�CG�;IG�;IP[GS�:RC��HfܷR66��R7g�R*V2��R&4��5@���U�H�NVDx�Du0�KF�LCTO���NN��OLw�ENuDY�LG;SLMx�FVRh�(�O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o�o�o�o# 5GYk}��� ������1�C� U�g�y���������ӏ ���	��-�?�Q�c� u���������ϟ�� ��)�;�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/�A�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� ������������ �'�9�K�]�o����� ������������# 5GYk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ����������%�1�STD~,�LANGM� H�`�r߄ߖߨߺ��� ������&�8�J�\� n����������� ���"�4�F�X�j�|� �������������� 0BTfx�� �����, >Pbt���� ���//(/:/L/�^$RBTL�OPT�Nu/�/�/�/�/�+DPNK��/�/??/? M�$�S?e?w?�?�?�? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q���������˟ݟ ���%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ����� /�A�S�e�wωϛϭ� ����������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy�� �����	- ?Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O__�99'U�$F�EAT_ADD �?	���TQ~\P  	$X e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������#�5GGTDEMO �RTY   $X������ ��///&/8/R/\/ �/�/�/�/�/�/�/�/ �/+?"?4?N?X?�?|? �?�?�?�?�?�?�?'O O0OJOTO�OxO�O�O �O�O�O�O�O#__,_ F_P_}_t_�_�_�_�_ �_�_�_oo(oBoLo yopo�o�o�o�o�o�o �o$>Hul ~������� � �:�D�q�h�z��� ����ݏԏ��
�� 6�@�m�d�v������� ٟП����2�<� i�`�r�������կ̯ ޯ���.�8�e�\� n�������ѿȿڿ� ���*�4�a�X�jϗ� �Ϡ����������� &�0�]�T�fߓߊߜ� �����������"�,� Y�P�b������� ��������(�U�L� ^��������������� �� $QHZ� ~�������  MDV�z� ������// I/@/R//v/�/�/�/ �/�/�/�/??E?<? N?{?r?�?�?�?�?�? �?�?
OOAO8OJOwO nO�O�O�O�O�O�O�O __=_4_F_s_j_|_ �_�_�_�_�_�_oo 9o0oBooofoxo�o�o �o�o�o�o�o5, >kbt���� ����1�(�:�g� ^�p�������ӏʏ܏ �� �-�$�6�c�Z�l� ������ϟƟ؟��� )� �2�_�V�h����� ��˯¯ԯ���%�� .�[�R�d�������ǿ ��п���!��*�W� N�`ύτϖ��Ϻ��� ������&�S�J�\� �߀ߒ߿߶������� ��"�O�F�X��|� ������������ �K�B�T���x����� ��������G >P}t���� ��C:L yp������ 	/ //?/6/H/u/l/ ~/�/�/�/�/�/?�/ ?;?2?D?q?h?z?�? �?�?�?�?O�?
O7O .O@OmOdOvO�O�O�O �O�O�O�O_3_*_<_ i_`_r_�_�_�_�_�_ �_�_o/o&o8oeo\o no�o�o�o�o�o�o�o �o+"4aXj� �������'� �0�]�T�f������� ��������#��,� Y�P�b����������� ������(�U�L� ^������������ܯ ���$�Q�H�Z��� ~��������ؿ�� � �M�D�Vσ�zό� �ϰ��������
�� I�@�R��v߈ߢ߬� ���������E�<� N�{�r�������� �����A�8�J�w� n������������� ��=4Fsj| ������ 90Bofx�� �����/5/,/ >/k/b/t/�/�/�/�/ �/�/�/?1?(?:?g? ^?p?�?�?�?�?�?�? �? O-O$O6OcOZOlO �O�O�O�O�O�O�O�O )_ _2___V_h_�_�_ �_�_�_�_�_�_%oo .o[oRodo~o�o�o�o �o�o�o�o!*W N`z����� ����&�S�J�\� v����������ڏ����"�O�F�r�  i��������� П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt����� ��(:L^>p  qk �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |������� ��0�B�T�f�x��� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� \�n������������� ����"4FXj |��������0BTfvzm����� ��/ /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo jo|o�o�o�o�o�o�o �o0BTfx �������� �,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vψ� �ϬϾ��������� *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx ������� ,>Pbt�� �����//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x���$FEAT_D�EMOIN  V{�����~���_INDEX��������ILECOM�P S����ޑ����ԐS�ETUP2 T�ޕ��  �N �ѓ_AP2�BCK 1Uޙ  �)y�G�V�%=�z�~��h��� {�<�ѯ`������+� ��O�ޯs������8� Ϳ߿n�ϒ�'�9�ȿ ]�쿁�ώϷ�F��� j���ߠ�5���Y�k� �Ϗ�߳���T���x� ���C���g��ߋ� ��,���P������� ��?�Q���u����(� ����^�����)�� M��q��6� �l�%�2[ ���D�h �/�3/�W/i/� �//�/@/�/�/v/? �//?A?�/e?�/�?�? *?�?N?�?�?�?O�?@=O�?JOsO�!�P%�� 2:�*.V1RzO�O2@*�O�O`/C�O_E�@PC_|H_2@FR6:3_"t^_�_'[T���_ �_]U�_�\���_o F�*.F�OOo1A	�_S=o|lo�o/kSTM�o�o\RbP�o }�o$/kH�oW�g�E�0jGIF ���e���-�0jJPG7�a��eM�
����(ZJS���2@�w�ҏ��%
Ja�vaScript�;�CS�h��fU��� %Casc�ading St�yle Shee�ts��@
ARGNAME.DTß
&L�`\ן�������ğ�DISP*���`[���*������H�
TPEIN�S.XML˯w�:�\߯����Cust�om Toolb�ar �O�PASS�WORD��$NF�RS:\c�"� %�Passwor�d Config ���?�|��#�YOG� ֿk�}�ϡ�0����� f��ϊ�߮���U��� y��r߯�>���b��� 	��-��Q�c��߇� ��:�L���p���� ��;���_������$� ��H�����~���7 ����m��� �� V�z!�E� i{
�.�Rd ��/�/S/�w/ /�/�/</�/`/�/? �/+?�/O?�/�/�?? �?8?�?�?n?O�?'O 9O�?]O�?�O�O"O�O FO�OjO|O_�O5_�O ._k_�O�__�_�_T_ �_x_oo�_Co�_go �_o�o,o�oPo�o�o �o�o?Q�ou ��:�^��� )��M��F������ 6�ˏݏl����%�7� Ə[���� ���D� ٟh�ҟ���3�W� i��������ïR�� v������A�Яe��� ^���*���N������ Ϩ�=�O�޿s�ϗ� &�8���\��π���'� ��K���o߁�ߥ�4� ����j��ߎ�#�����Y�;��$FILE�_DGBCK 1�U��F���� < ��)
SUMMAR�Y.DGc��M�D:�����D�iag Summ�ary����
CONSLOG�������[���Console log\����	TPACCN�Q���%������T�P Accoun�tin}���FR�6:IPKDMPO.ZIP�
'�`����Excep�tiond��MEMCHECK���8����o�Mem�ory Data��;�YF)	FTPN�?�C��q�mment �TBDl;�L =��)ETHERNETa������Ethern�et s�figu�ra���VDCSVRF`FXq/��%6  verify allt/�>�M+�1%DI�FFi/O/a/�/� {%�(diff�/��'�6 CHG01 �/�/�/{?�!?�?�"*f992q?X?j?�?
?�?�?@23�?�?�?��O O�O9F�VTRNDIAG.LS�O`OrO_���A ��nost�ic_>�T6a�)UPDATE�S.MP3_�FR�S:\K_�]��U�pdates L�ist�_�PSRBWLD.CM�_��wR�_�_p�PS�_ROBOWEL����AHADO�W�O�O�O�o�S�hadow Ch�anges�o{qQbNOTI;/�lo~o�Not�ific"�o;�+@AG��j�9� �����w��� B��f�x����+��� ҏa��������'�P� ߏt������9�Ο]� ����(���L�^�� �����5���ܯk� � ��$�6�ůZ��~��� ���C�ؿ�y�ϝ� 2���?�h�����ϰ� ��Q���u�
�߫�@� ��d�v�ߚ�)߾�M� ���߃���<�N��� r����7���[��� ���&���J���W��� ���3�����i����� "4��X��|� �A�e��0 �Tf���� O�s//�>/� b/�o/�/'/�/K/�/ �/�/?�/:?L?�/p? �/�?�?5?�?Y?�?}? �?$O�?HO�?lO~OO �O1O�O�OgO�O�O _ 2_�OV_�Oz_	_�_�_ ?_�_c_�_
o�_.o�_ Rodo�_�oo�o�oMo �oqo�o<�o` �o��%�I�� ��8�J��n�� ��!���ȏW��{�� "���F�Տj�|���� /�ğ֟e�������� +�T��x������=� үa������,���P� b�񯆿���9���� o�ϓ�(�:�ɿ^�� �ϔ�#ϸ�G�����}πߡ�6���C�l�N���$FILE_FR�SPRT  ���V�������MDONL�Y 1U��N�� 
 �)MD�:_VDAEXTP.ZZZs�$����
�6%NO� Back fi�le ��N�S�6�\��߀�Iߍ�� ����i������4��� X�j���������S� ��w���B��f ����+�O�� ��>P�t �'��]��/ (/�L/�p/�//�/�5/�/�/��VISB�CK�؝���*.�VD�/'?� FR�:\� ION\DOATA\?�"� �Vision VD(�S?a/�?�?�/ �?�/�?�?O+O�?OO �?sO�OO�O8O�O\O nO_�O'_9_�O]_�O �__�_�_F_�_j_�_ o�_5o�_Yo�_�_�o o�o�o�o�oxo�o C�og�o��,��P�t��{�L�UI_CONFIoG V��	1>&� $ ���{��}�������ŏ׏�e�|x��!�3� E�W�g����������� ҟi����,�>�P� �t���������ίe� ���(�:�L��p� ��������ʿa�� � �$�6�H�߿l�~ϐ� �ϴ���]������ � 2�D���h�zߌߞ߰� ��Y�����
��.��� ?�d�v����C��� ������*���N�`� r�������?������� &��J\n� ��;���� "�FXj|�� 7����//� B/T/f/x/�/!/�/�/ �/�/�/?�/,?>?P? b?t?�??�?�?�?�? �?O�?(O:OLO^OpO �OO�O�O�O�O�O _ �O$_6_H_Z_l_~__ �_�_�_�_�_�_�_ o 2oDoVohozoo�o�o �o�o�o}o�o.@ Rd�o����� �y��*�<�N�`� ���������̏ޏu� ��&�8�J�\�󏀟 ������ȟڟq���� "�4�F�X��|�����в�į֯f��|��$FLUI_DA�TA W��}��j����RESULT �2X�0� ��T�/wiz�ard/guid�ed/steps/Expert� g�y���������ӿ����	��)��Co�ntinue w�ith GD�ance)�d�vψϚϬπ����������*� ��-��I�0 �r�I�	��i��;�ps,ߴ��� ������� �2�D�V� h�z�9�r�������� ������1�C�U�g�@y���i�[�m����torch�� %7I[m�� ������!3 EWi{���������������wproc��U/g/y/�/ �/�/�/�/�/�/	?? �??Q?c?u?�?�?�? �?�?�?�?OO)O���DO/����M�T�imeUS/DST3O�O�O�O�O__�'_9_K_]_o_2�DisablRϤ_�_ �_�_�_�_o"o4oFo�Xojo|n�j��eOWOiO{O�O�B24 �O/ASew ����~_�_�� �+�=�O�a�s����� ����͏�o�o�o�o���:�L�Region Џ_�q���������˟�ݟ���.�AmericaI/M�_� q���������˯ݯ���.�ہyE���]�8�1��BEdi��$� ��ſ׿�����1��C�U�g�*; Tou�ch Panel� �� (reco/mmen��)uϺ� ��������&�8�J�\�n�-��=�O���s�|���Bacces<� ��*�<�N�`�r������)<Con�nect to Network��  ��$�6�H�Z�l�~� ��������1��鏣�����!�ߝ@IntroductK� ^p������ � -?6HZl ~�������/ / =O��=/ �b0�/�/�/�/�/�/ �/?#?5?G?Y?k?* �?�?�?�?�?�?�?O@O1OCOUOgO׈@ |]/G*���~�O �O}/�O�O__*_<_ N_`_r_�_�_�_�_y? �_�_oo&o8oJo\o no�o�o�o�ouO�O�O �O�O4FXj| �������� �_0�B�T�f�x����� ����ҏ������o �o�o_�!�������� Ο�����(�:�L� ^����������ʯܯ � ��$�6�H�Z�l� +�=�O���s�ؿ��� � �2�D�V�h�zό� �ϰ�o�������
�� .�@�R�d�v߈ߚ߬� ��}��ߡ��ſ*�<� N�`�r������� ������%�8�J�\� n��������������� ����1��U�| ������� 0BTf%��� �����//,/ >/P/b/!�/E�/i k/�/�/??(?:?L? ^?p?�?�?�?�?w�? �? OO$O6OHOZOlO ~O�O�O�Os/�O�/�O _�?2_D_V_h_z_�_ �_�_�_�_�_�_
o�? .o@oRodovo�o�o�o �o�o�o�o�O_�O 3]_����� ����&�8�J�\� o��������ȏڏ� ���"�4�F�X�a ;����q֟���� �0�B�T�f�x����� ��m�ү�����,� >�P�b�t�������i� {������ß(�:�L� ^�pςϔϦϸ����� �� ߿�$�6�H�Z�l� ~ߐߢߴ��������� �Ϳ߿�S��z�� �����������
�� .�@�R��v������� ��������*< N`�1�C�g�� ��&8J\ n���c���� �/"/4/F/X/j/|/ �/�/�/q�/��/� ?0?B?T?f?x?�?�? �?�?�?�?�?O?,O >OPObOtO�O�O�O�O �O�O�O_�/%_�/I_ ?p_�_�_�_�_�_�_ �_ oo$o6oHoZoO ~o�o�o�o�o�o�o�o  2DV_w9_ �]__���
�� .�@�R�d�v������� koЏ����*�<� N�`�r�������gɟ ����Ï&�8�J�\� n���������ȯگ� ����"�4�F�X�j�|� ������Ŀֿ����� �ݟ'�Q��xϊϜ� ������������,� >�P��t߆ߘߪ߼� ��������(�:�L� �U�/�y��e����� �� ��$�6�H�Z�l� ~�����a���������  2DVhz� �]�o������ .@Rdv��� ������/*/</ N/`/r/�/�/�/�/�/ �/�/?���G?	 n?�?�?�?�?�?�?�? �?O"O4OFO/jO|O �O�O�O�O�O�O�O_ _0_B_T_?%?7?�_ [?�_�_�_�_oo,o >oPoboto�o�oWO�o �o�o�o(:L ^p���e_��_ ��_�$�6�H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ����� �=��d�v������� ��Я�����*�<� N��r���������̿ ޿���&�8�J�	� k�-���Q�S������� ���"�4�F�X�j�|� �ߠ�_���������� �0�B�T�f�x��� [Ͻ��������,� >�P�b�t��������� ��������(:L ^p������ �������E�l ~������� / /2/D/h/z/�/ �/�/�/�/�/�/
?? .?@?�I#m?�?Y �?�?�?�?OO*O<O NO`OrO�O�OU/�O�O �O�O__&_8_J_\_ n_�_�_Q?c?u?�?�_ �?o"o4oFoXojo|o �o�o�o�o�o�o�O 0BTfx�� ������_�_�_ ;��_b�t��������� Ώ�����(�:��o ^�p���������ʟܟ � ��$�6�H��� +���O���Ưد��� � �2�D�V�h�z��� K���¿Կ���
�� .�@�R�d�vψϚ�Y� ��}��ϡ���*�<� N�`�r߄ߖߨߺ��� ������&�8�J�\� n����������� �����1���X�j�|� �������������� 0B�fx�� �����, >��_!��E�G� ���//(/:/L/ ^/p/�/�/S�/�/�/ �/ ??$?6?H?Z?l? ~?�?O�?s�?�?�/ O O2ODOVOhOzO�O �O�O�O�O�O�/
__ ._@_R_d_v_�_�_�_ �_�_�_�?�?�?o9o �?`oro�o�o�o�o�o �o�o&8�O\ n������� ��"�4��_=ooa� ��Mo��ď֏���� �0�B�T�f�x���I ����ҟ�����,� >�P�b�t���E�W�i� {�ݯ����(�:�L� ^�p���������ʿܿ �� ��$�6�H�Z�l� ~ϐϢϴ������ϩ� ��ͯ/��V�h�zߌ� �߰���������
�� .��R�d�v���� ����������*�<� ���߁�Cߨ����� ����&8J\ n�?����� �"4FXj| �M��q�����/ /0/B/T/f/x/�/�/ �/�/�/�/�??,? >?P?b?t?�?�?�?�? �?�?�O�%O�LO ^OpO�O�O�O�O�O�O �O __$_6_�/Z_l_ ~_�_�_�_�_�_�_�_ o o2o�?SoOwo9O ;o�o�o�o�o�o
 .@Rdv�G_� ������*�<� N�`�r���Co��goɏ ۏ���&�8�J�\� n���������ȟڟ� ���"�4�F�X�j�|� ������į֯��ߏ�� �-��T�f�x����� ����ҿ�����,� �P�b�tφϘϪϼ� ��������(��1� �U��A��߸����� �� ��$�6�H�Z�l� ~�=Ϣ���������� � �2�D�V�h�z�9� K�]�o�������
 .@Rdv��� �����*< N`r����� �������#/��J/\/ n/�/�/�/�/�/�/�/ �/?"?�F?X?j?|? �?�?�?�?�?�?�?O O0O�//uO7/�O �O�O�O�O�O__,_ >_P_b_t_3?�_�_�_ �_�_�_oo(o:oLo ^opo�oAO�oeO�o�O �o $6HZl ~������o� � �2�D�V�h�z��� ����ԏ�o���o� �o@�R�d�v������� ��П�����*�� N�`�r���������̯ ޯ���&��G�	� k�-�/�����ȿڿ� ���"�4�F�X�j�|� ;��ϲ���������� �0�B�T�f�x�7��� [����ߓ�����,� >�P�b�t����� �������(�:�L� ^�p������������� �߭���!��HZl ~�������  ��DVhz� ������
// ��%��I/s/5�/�/ �/�/�/�/??*?<? N?`?r?1�?�?�?�? �?�?OO&O8OJO\O nO-/?/Q/c/�O�/�O �O_"_4_F_X_j_|_ �_�_�_�_�?�_�_o o0oBoTofoxo�o�o �o�o�o�O�O�O�O >Pbt���� ������_:�L� ^�p���������ʏ܏ � ��$��o�oi� +������Ɵ؟��� � �2�D�V�h�'�y� ����¯ԯ���
�� .�@�R�d�v�5���Y� ��}������*�<� N�`�rτϖϨϺ��� ݿ����&�8�J�\� n߀ߒߤ߶��߇��� ���Ͽ4�F�X�j�|� ������������� ���B�T�f�x����� ������������ ;��_!�#��� ���(:L ^p/������ � //$/6/H/Z/l/ +�/O�/�/��/�/ ? ?2?D?V?h?z?�? �?�?�?��?�?
OO .O@OROdOvO�O�O�O �O}/�/�/�O_�/<_ N_`_r_�_�_�_�_�_ �_�_oo�?8oJo\o no�o�o�o�o�o�o�o �o�O_�O=g)_ �������� �0�B�T�f�%o���� ����ҏ�����,� >�P�b�!3EW�� {�����(�:�L� ^�p���������w�ܯ � ��$�6�H�Z�l� ~�������ƿ������ �͟2�D�V�h�zό� �ϰ���������
�ɯ .�@�R�d�v߈ߚ߬� ����������׿� ��]�τ������ ������&�8�J�\� �m������������� ��"4FXj)� �M�q���� 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ {�/�?�(?:?L? ^?p?�?�?�?�?�?�? �? OO�6OHOZOlO ~O�O�O�O�O�O�O�O _�//_�/S_?_�_ �_�_�_�_�_�_
oo .o@oRodo#O�o�o�o �o�o�o�o*< N`_�C_��{o ����&�8�J�\� n���������uoڏ� ���"�4�F�X�j�|� ������q��ߟ	� �0�B�T�f�x����� ����ү����Ǐ,� >�P�b�t��������� ο���ß��1� [���ϔϦϸ����� �� ��$�6�H�Z�� ~ߐߢߴ��������� � �2�D�V��'�9� Kϭ�o�������
�� .�@�R�d�v������� k�������*< N`r����y� ������&8J\ n������� ���"/4/F/X/j/|/ �/�/�/�/�/�/�/? ���Q?x?�?�? �?�?�?�?�?OO,O >OPO/aO�O�O�O�O �O�O�O__(_:_L_ ^_?_A?�_e?�_�_ �_ oo$o6oHoZolo ~o�o�o�o�_�o�o�o  2DVhz� ��o_��_��_� .�@�R�d�v������� ��Џ����o*�<� N�`�r���������̟ ޟ���#��G�	� ���������ȯگ� ���"�4�F�X��|� ������Ŀֿ���� �0�B�T��u�7��� ��o���������,� >�P�b�t߆ߘߪ�i� ��������(�:�L� ^�p����eϯω� �����$�6�H�Z�l� ~��������������� �� 2DVhz� ��������� ��%O�v��� ����//*/</ N/r/�/�/�/�/�/ �/�/??&?8?J?	 -?�?c�?�?�? �?O"O4OFOXOjO|O �O�O_/�O�O�O�O_ _0_B_T_f_x_�_�_ �_m??�?�_�?o,o >oPoboto�o�o�o�o �o�o�o�O(:L ^p������ � ��_�_�_E�ol� ~�������Ə؏��� � �2�D�U�z��� ����ԟ���
�� .�@�R��s�5���Y� ��Я�����*�<� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ�c��χ��� ���"�4�F�X�j�|� �ߠ߲��������߹� �0�B�T�f�x��� �������������� ;�����t��������� ������(:L �p������ � $6H�i +���c���� / /2/D/V/h/z/�/ �/]�/�/�/�/
?? .?@?R?d?v?�?�?Y �}�?�?�O*O<O NO`OrO�O�O�O�O�O �O�O�/_&_8_J_\_ n_�_�_�_�_�_�_�_ �?�?�?oCoOjo|o �o�o�o�o�o�o�o 0B_fx�� �������,� >��_o!o3o��Wo�� Ώ�����(�:�L� ^�p�����S��ʟܟ � ��$�6�H�Z�l� ~�����a�s���篩� � �2�D�V�h�z��� ����¿Կ濥�
�� .�@�R�d�vψϚϬ� �������ϳ�ůׯ9� ��`�r߄ߖߨߺ��� ������&�8���I� n����������� ���"�4�F��g�)� ��M߲��������� 0BTfx�� ������, >Pbt��W�� {����//(/:/L/ ^/p/�/�/�/�/�/�/ �/�?$?6?H?Z?l? ~?�?�?�?�?�?�?� O�/O��?hOzO�O �O�O�O�O�O�O
__ ._@_�/d_v_�_�_�_ �_�_�_�_oo*o<o �?]oO�o�oW_�o�o �o�o&8J\ n��Q_���� ��"�4�F�X�j�|� ��Mo�oqo��叧o� �0�B�T�f�x����� ����ҟ䟣��,� >�P�b�t��������� ί௟��Ï�7��� ^�p���������ʿܿ � ��$�6���Z�l� ~ϐϢϴ��������� � �2����'��� K�����������
�� .�@�R�d�v��GϬ� ����������*�<� N�`�r�����U�g�y� ����&8J\ n�������� �"4FXj| ���������� ��-/��T/f/x/�/�/ �/�/�/�/�/??,? �=?b?t?�?�?�?�? �?�?�?OO(O:O� [O/OA/�O�O�O�O �O __$_6_H_Z_l_ ~_�_�O�_�_�_�_�_ o o2oDoVohozo�o KO�ooO�o�O�o
 .@Rdv��� ����_��*�<� N�`�r���������̏ ޏ�o���o#��o�\� n���������ȟڟ� ���"�4��X�j�|� ������į֯���� �0��Q��u���K� ����ҿ�����,� >�P�b�tφ�E��ϼ� ��������(�:�L� ^�p߂�A���e����� �� ��$�6�H�Z�l� ~����������� � �2�D�V�h�z��� �����������߷� +��Rdv��� ����*�� N`r����� ��//&/����	 }/?�/�/�/�/�/ �/?"?4?F?X?j?|? ;�?�?�?�?�?�?O O0OBOTOfOxO�OI/ [/m/�O�/�O__,_ >_P_b_t_�_�_�_�_ �_�?�_oo(o:oLo ^opo�o�o�o�o�o�o �O�O�O!�OHZl ~������� � ��_1�V�h�z��� ����ԏ���
�� .��oO�s�5���� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���?���c�ſ��� ���"�4�F�X�j�|� �Ϡϲ����ϕ���� �0�B�T�f�xߊߜ� �����ߑ��ߵ��ٿ ��P�b�t����� ��������(���L� ^�p������������� �� $��E�i {?�������  2DVhz9� ������
// ./@/R/d/v/5Y �/�/��/??*?<? N?`?r?�?�?�?�?�? ��?OO&O8OJO\O nO�O�O�O�O�O�/�/�/�O_%Q�$FM�R2_GRP 1�Y%U� ��C4  B]��0	 �0c_�u\`PF�6 F@�S�Q�T�J`S�_�]�`P?�  �_�_<�P�a;O��O9 n�e�]A`l+o=kBH]SB�YP<X`;a@�33ce�\��_�o�Y@UO� �a�o�_�o�o�o�o 4XC|g�����}9R_CFG {ZF[T ���(�:��{NO �FZ
F0p� �u��|RM_CHK?TYP  6Q�0pNPPPP8QROM���_MIN���3������|`X9PSS�B�s[%U aV��5�
����uTP_DEF�_OW  �4|NS1�IRCOM���B��$GENOV_RD_DO���1no�THR�� d���du�_ENBa� �u�RAVC?S\:Ӈހ ��U"���1��?�P�sj� �ՑOUBPb�F\x�sXF�sU<�� �]ǯq�������3C�YP��YP�%��d��1A@M�?�U�vY��#�֐SMT?Sc�RP���4��$HOSTC��r1dFY߀���? 	
�
�d
��6:��9eV� �ϙϫϽ���u��� ���$�G�H���	anonymousK� yߋߝ߯��� 	�� -�
�A�c���R�d�v� ���Ϭ��������� M�_�<�N�`�r����� ��������7�& 8J\����� ���!�3�"4F X��������� ��//e//T/f/ x/�/��/��/�/�/ ??as���/s? ��?�?�?�?�?9/O (O:OLO^O�?�/�/�O �O�O�O�O5?G?Y?_ mOZ_�?~_�_�_�_�_ q_�_�_o oC_Do�O hozo�o�o�o�O	__ -_
Aoc_@Rdv ��_����� Mo_o<�N�`�r����o �o�o���7�&� 8�J�\���������� ُǟ!����"�4�F�����ENT 1e��� P!ڟ��  ����ï��� ���ί/��;��d� ��L���p�ѿ������ �ܿ�O��s�6ϗ� Zϻ�~ϐ��ϴ���� 9���]� �Vߓ߂߷� z��ߞ��������4� Y��}�@��d���� �������C��g��*�QUICC0 t�P�b�����1��������2��c�!ROUTER�d@R�!PC�JOG��!�192.168.�0.10����CA�MPRT�!b�1� +RT}�/A�h�NAME� !u�!RO�BO�S_CF�G 1du� ��Auto�-started^��FTP��;! ͏ϟf/��/�/�/�/ �/o��/??,?O/=? �/t?�?�?�?�?��/ &/8/OL?n/,O]OoO �O�OZ?�O�O�O�O�O "O�O5_G_Y_k_}_�_ ������ʏ_�_BOo 1oCoUogo._�o�o�o �o�o�_xo	-? Qc�_�_�_��o� o���)��oM�_� q������:���ݏ� ��%�l~���� �����ǟٟ���ď !�3�E�W�i������ ��ïկ���@�R�d� A�x�e����������� ��|�����+�N�O� �sυϗϩϻ��� &�8�:��n�K�]�o� �ߓ�ZϷ��������� "ߤ�5�G�Y�k�}�� �����Ϩ����B�� 1�C�U�g�.������ ������x�	-?�Q��_ERR �f�aqPDU�SIZ  ��^����>�WR�D ?%��� � guest����)�;�SCD_GR�OUP 3g, u!�� ��LOA��RE�S�TM� $v�T_�ENBs �TTP_AUTH� 1h� <!�iPendan�GR.���A!KAREL:*R/[/m-KC�/�/�/�z VISION SETk?�/F!??1?w#U?C?m? g?�?�?�?�?�?�>!$CTRL i��;H��
��F�FF9E3�?���FRS:DEFA�ULT`LFA�NUC Web ?Server`JNB !$��	L�O�O�O_�_,_oWR_CONFIG jp��`OqI�DL_CPU_P5C@��B����Pw BH�UMIN�\�x�UGNR_IO�z�����PNPT_SIM_DO�V��[STAL_S7CRN�V �6F�Q�TPMODNTOqLg�[�ARTY�X@�Q�V� %  gx��SOLNK 1k�}�o�o�o�o�o� �bMASTE��Pzi�UOSLA�VE l�AuRAMCACHE0�(bO'!O_CFGr�c�sUO0��r�CYCLq�uy@_?ASG 1maW�
 �)�;�M� _�q���������ˏݏp��{�rNUM�5�	
�rIPo�wRTRY_CN@��R�
�ra_UPD��a�� �r�p�r�nP~u��u�PS�DT_ISOLC�  P{v"�J_23_DSrd.N��OGg1oP{�<��d<�P� #?��R��?�����Q��̯ޯ𯯯�&�8�J�������*�ЮP�qi��PhpEC�so�UKANJI_�*pK�_³� MONG pp;_��y� (�:�L�^�pϒ~"���qa\EF�ŭ���C�L_L�P'�J�İEYLOGGIN�p�u�F���$�LANGUAGE� �FabyD l<�qLG�qr�y^�a ���xu ��e����P���'U0�����;��cM�CH ;��
��(?UT1:\���� ���������!�@3�E�\�i�{��(����lLN_DISP sP�ئ���f��OC4b�RDz�S��A@�OGBOO/K tM�d��>A���k�X�܏��� ������<O�Y���	>F	Q������N�`��O�_BUFoF 1u�me2kE�j�FB�iG� �G>P} t������/�//C/��~DCS� w�{�=���G��/�/�/|�/Z$IO 1x�{G ğ3D��? *?<?N?b?r?�?�?�? �?�?�?�?OO&O:O JO\OnO�O�O�O�O�OZ�%E�PTM�dh� #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo1o�CoUogoyo�o-��BS�EV�����FTYP�_�o�m���RSh���|��F�L 2y=��� �/�������F(TP����b'�NGNAM�6%.�nV$UPS��GIh������f�_LOA�DPROG %���%	T_ARC�WEL�����MA?XUALRM'��A85�̀l�_PRh���� E�	ˀC��z�M�������,�P �2{� ت	Z�aڀ	�|�f4� �~����������(Ο ���3��(�i�T��� x���ï���ү��  �A�,�e�P�����~� �����ƿؿ��=� (�a�s�VϗςϻϞ� ������� �9�K�.� o�Zߓ�v߈��ߴ��� ���#��G�2�k�N� `������������ �
�C�&�8�y�d��� ������������ć�DBGDEF �|$�:!"�$6 _L?DXDISAQ�#���#MEMO_AP�K�E ?$�
 H�������"ˀISCW 1}$�%�� oy�M�����QE_MSTR �~�m%SCD 1���T/�x/ c/�/�/�/�/�/�/�/ ??>?)?b?M?r?�? �?�?�?�?�?O�?(O O%O^OIO�OmO�O�O �O�O�O _�O$__H_ 3_l_W_�_{_�_�_�_ �_�_o�_2ooBoho So�owo�o�o�o�o�o �o�o.R=va ����������<�'�`��MJPTCFG 1�+�]�%�����MI/R 1�%Ԁp�@T�q���T��< G ?� �%��t�7�q�� i������������� 1�C�֟��j�L�V�x� ��P�����ί��0� T�E �q����8��� ������򿐿����  �B�p�R��ϵ���Z� |���п����6���>� l�R�d߆߈ߖ����� �ߞ���2���@�z� `����������� +�=��������X�b� t�������������* ��o�6��� ������
 @nP���Xz ����4/�,/j/@P/b/�/�/���K��;���  �/���LTARM_�"�̅� �"����6?�>4��METPU ; T����%���NDSP_ADC�OLX5� c>CMN�Ty? l5MST ��-�?���!�?|�4l5POSCF�7=�>PRPM�?�9[STw01���4܁<#�
gA[�gEwO �GcO�O�O�O�O�O�O _�O_G_)_;_}___�q_�_�_�_�_�Ql1S�ING_CHK � |?$MODAQ3����,�.#e�DEV 	��	�MC:WlHSI�ZEX0�-�#eTA�SK %��%$�12345678�9 �o�e!gTRI������ l̅% &�O2}���c�YP�a��9d"cE�M_INF 1��7;a`)AT&FV0E0X��})�qE0V1�&A3&B1&D�2&S0&C1S�0=�})ATZ�#�
�H'�O��qCw��A���b�ˏ���� �&���� ���3���ۏȟڟ�� ����"�4��X��� ��A�S�e�֯៛�� C�0����f�!���q� ����s�俗�����ͯ >��bϙ�sϘ�K��� w��������ɿۿL� ���#ϔߦ�Y���� �ߩ߳�$���H�/�l� ~�1ߢ�U�g�yߋ��� �� �2�i�V�	�z�5����������PoNIT�OR�0G ?kk �  	EXESC1�223E45�`789�� �(�4�@� L�X�d�p�T|�2�2�2�U2�2�2�2�U2�2�2�3��3�3(#aR_G�RP_SV 1��{ (�Q����<�qI�?b��@H|?�u��@4]$Rm�a_�Ds�n�ION_�DB-`�1m�1 � �K`�Fh"%B�++��0.Fh��N� Bl"$ Fi-ud1}e�/�/�/1�PL_NAME �!�e� �!�Default �Personal�ity (fro�m FD)b"P0R�R2� 1�L?68L@P�!K`
 d�2-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO�O�O�Of#2)?�O�O �O__,_>_P_b_t_f"<�O�_�_�_�_�_ �_
oo.o@oRodotl&�" �_�n
�o�of$P�o�o $6 HZl~���� ����o�o2�D�V� h�z�������ԏ� ��
��.�@��!�v� ��������П���� �*�<�N�`�r�����1e����ïխf"d��������(� 6����� �m���j���V� ������Ŀ ֿ�����:Ϸ�]�4m�f"��	`��������σ�:�oA�b)�����c' �A�  /�	23���)X ���E� ��X�, @D�  &t�?�z�n�?f |�f!AI�t�j���;�	l��	 �� � �h�Y Z ����� � x? � � ��ҷ�K_K }�K7X�K���J��?J�+����%��ԯC�@��6@�
�\��?(E@�Sє���.��=�N��������T;f�a�����$���*  ´  ��1�>�����z�w����<�
���� �Z!/���1�y�D�  �  ��  �`�#�H �l����-�	'�� � ��I�� �  ��0�&�:�È��ß�=�����0�@����%�f����f�(�2�+�a!v � '�Y��@!�p@���@��@��@��C��C�� �� C��C���C��f ��A���=����u"T�Bb $/��Lf!Dz��o��~�@��������A �л�D�  X ,>f �?�ffG�*/</� }�q/�+1��8~`�/�*>��H$��(�(~`�%P�(�������>�$����W�<�	<S��;�9<���<#*o<���M,@�K;|���f��",�?fff�? ?&�0T�@��.�2�J<?N\��55	��1��(� |��?z��?j7��[/0O OTO?OxOcO�O�O�O`�O�O�O{h�5F�� �O2_�OV_�?w_�9I_ �_E_�_�_�_�_oo oLo7opo[o�oo�o �oU�o�o��m_3�_�Z�o~���O*��& Q/�wl��q
��m.��+�d�V���Aa0��5uCP���L�<č?�����#��Y�/Ӄj6�B]�D��CC3�� z���������@I��l����A���A��PA ��R?�1>��-8��������O\����Q����#�
؞���A�иRA���C;���Q섟�"\)C0����qBo
=���Q�����8�Hp��G�� H�0�H��E1� C�&��Hy��I���H��%F�� �E,�s�]�i�E�I��@H����H��E# D�7�د�կ� ��2��V�A�z�e�w� ����Կ������� @�R�=�v�aϚυϾ� ����������<�'� `�K߄�oߨߺߥ��� �����&��J�5�G� ��k���������� �"��F�1�j�U��� y������������� 0T?x�u� �����tP�(�3�(���	4���<�̷�t�Ӂ3���8����ʭ���Ӂ� &n�
/4�f4yϱ$- $)d/R/�/v/�/�,Յ%PD2P�.�a�o?@Z?=?(?a?L<?g?�n?�?�?�?�?�?  �����?�?+OO OO:OsO?�o�O�O�O�L7�O�O_�O _F_4_JQ�L_^_�_�_p�_�_�_�Z  2jO�o  B��}���Cq���Ӏ@��RoӀ�Mqko}o�o^o�oҌ o�o�o/Aӄ��TӀӀ�a:Ӏ؎
 I� �������)��;�M�_�q����sq ����1��"��$MSKCFMA�P  $%� �Vsqoq����ONREL  ��%Ӂ�P��E�XCFENB�
у���FNy�'���JOGOVLIM��d��d��KE�Y�q�z�_P�AN�������RU�Na���SFSP�DTY� '����S�IGN��T1M�OTc����_C�E_GRP 1�$%Ӄ\dOh�\O �����T��ɯ���� �#�گG���<�}�4� ����j�׿�����Ŀ 1��*�g�ϋϝτ� ��x���������f��QZ_EDIT��͇��TCOM_C_FG 1�ɍ~v�v߈ߚ�
V�_AR�C_"��%P�T_MN_MODE���0�UAP_C�PL��4�NOCH�ECK ?ɋ �%�3�E�W� i�{���������������/�A��NO_WAIT_L�lK�6�NT^��ɋ�u|��_ERR@�29�ɉ�Q� ��������4F���MO����|t5����*�XEB���C3�B�ƀC!xX�<���?�l�K�np����PARAM���ɋ�/`�2t8�_^ =�P�345678901x��s��� �//�9/K/'+t7��}/�,"�/��ODRDSP���0��OFFSET_C�ARA���&DIS��/�#S_A��AR�K�L�OPEN_FILE0h���L����OPTION_�IO����m0M_P�RG %Ɋ%$�*�?�>I3WO50-�F�0� �5D���2��0@�'A	 ���C���#��� RG_DS�BL  Ʌ��v|rO�!RIENTkTO��!C�mp�ҁ,a� UT_SIM_Du7Ђ��� �V� LCT � ��H��4���I�%y��A�_PEX��?TR[AT�� d0�T>� UP ��N�pK��i_{_XrfS`�bgq�Rn�}]�$��2?��L68L�@P�C
 d�/�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\��2�_������ �
��.��{X�j� |�������ď֏��� ����H�X��PX�~��"Pk�����̟ޟ ���&�8�J�\�n� ��������������� �"�4�F�X�j�|��� ����Ŀֿ���ɯۯ 0�B�T�f�xϊϜϮ� ����������,�>���E�}ߏ�SI�߿ޤ�����b�@bݢ/3��W�
�@ L�v�l�~��������J�Q�'�)L�	�``�Z�l�~���:�o�A��������KA�  ���T�P�OOP1�[��v��TH��E=D�X, @D� � 2��,?�D�4429�h;�	�l�	@� �� �h��_`� �� �� x � � ���JH�H�2�-HL��H��lH�WG���=�3Ho���JC��@p�@ע�@�P1���0�Z�@�S �>PP@%ICUB��<� �K��@��a��y�  ��  �  �
 #�0�*&�H/�	'� � f"�I� �  �����=���8�/�+�@�/�  �>A�/M+>B��r�N�@4?  'x0�L4�0C�@C��+ CC�C�Y?�k?D�  �A��!����~����B�@�1�����!
ENz�-O�QO<OaO�O�^/p(�1�E�S� ��<��1�P.   �?�ff��O�O�OC 7�/_A[sA8��W_eZ>�' �$FjJ(��UP�X�I@����#�T[���<�	<S��;�9<��<#*o<��5��\@�	k:���#�R��?fff?�� ?&D`�@�.�Vb�J<?N\�be:��2?aKjI: �o8�o(g~_�o�o �o6!ZE~� {�������o �o�o�h����w��� ��ԏ��я
���.�� R�=�v�a�?��o�e +��O����<�N�`��r�Z���@_��l � /�ȯ+��ׯ�"�����A`>��?�C��s�
�П��?��ء����̿n	�/VX���B�D90#CC�ޚ��������^�@I�*�����A��A���PA �R?��1>�-�������ÍO\����Q����#�
������AиRA����C;����Q�B��0\)C�0���qB�o
=��Q�������Hp���G� H�0��H��E1� �C���Hy��I���H��%F?�� E,�1߯�i�EI��@H����H��E?# D����� �ߓ��߷�������� 8�#�5�n�Y��}�� �����������4�� X�C�|�g��������� ������	B-f xc������ �>)bM� q�����/� (//L/7/p/[/m/�/ �/�/�/�/�/?�/6? H?3?l?W?�?{?�?�?��?�?�?O��(��33�([��T��BE�5��̷�2ODOX�3ǲ��^OpO~B���O�OX�� &n��O�O4�f4yϱ�M�I"__F_4_(j_X\��PbP�^�����_O�_�_�_o
l?%o,oeoPouo�o~�o  ���ʞo �o�o�o�o1�_��dR�v|7���`�������
���R�@�v�d����� s 2(я  BG��;�G�C/�D�X�@ K��"�4�F�X�j�{���������ɟ۟�T��X���X�X�ꕑX���
  �W�i�{�������ï կ�����/�A����1� ���K1���"�$PARAM�_MENU ?��E� � MNUT�OOLNUM[1-]݆��F~������AWEPC�R��.$INCH�_RATE��S�HELL_CFG�.$JOB_BA�S߰ WVW�PR.$CENTER_RI�������AZIMUTH �OPTB����E�LEVATION� TC����DW��TYPE SN��ARCLINK�_AT �STAT�USǳ]�__VA�LU߱̰LEP>��.$WP_���� �U�̢ϴ��������π�7�2�D�V��z�S�SREL_ID � �E�Q���US�E_PROG �%��%{��ߏ�CC�RT�ԶQ����_H�OST !��!��5���T�P��Q���*�S����_T�IMEOU�Ս� � z�GDEBU�G�Љ���GINP?_FLMSK����TR����PGd� e ����$�CH��(��Q���z�t� ����������( :c^p���� ��� ;6H Z�~�������// /2/[/��W�ORD ?	��
? 	RS�C�PNn�BMA�IW��#SU&��#T�Et�CSTYL COL0eW(�/�W�TRACECToL 1��E��� �P�P7D/T Q��ED0!0�D � �S���QQ6� [;q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ� ���#�5�G�Y�k�}��6LEW���5���3  �6_UPg �<;b������ ���&�0��M$a��R�\0R� � ��)_DEF�SPD ���2���  �z�I�NؐTRL ����a�8!�h�PE__CONFIܐ�7����M!b,L�IDٓ���	ĨG�RP 1�9 �lM!A>ff���\�
=�D�  DZ� kD
�@�
�M �d!�?�O��������H�"�$�i� ´����m�B��̱����ਿ�̿��&�B34�$�]�o�Y� <<j��tϭ� pϪ�������ό��@O��_߅�p��z����M 
���ߊ���� ��5� �Y�D�}�h�� ������������*��)<�
V7.1�0beta1��� A�k�\�B�
��(�Y�?&f�fp�>.{X��
�����X�B!�념�A{33A�&�(�h� -������������pM"�Ȁ3EWM$ғ�K�NOW_M  �0��ȤSV �.:�%��� ����IM"TG��M�=�(��	������.�* ��ś�M#�)�Y�@ )���M % .ѐȡMR�=�$��հ�f/x+��ST�1� 1�<9^ 4 �()�o��/�/�/
? �/?!?S?E?W?�?{? �?�?�?�?O�?�?>O�O/OtOSOeOwO�'2p�,��/���<�O�O� 3�O�O�O�O�'A4_-_?_Q_�'5n_�_�_�_�'6�_�_�_�_�'7o&o8oJo�'�8goyo�o�o�'MA�D�� ȕ�EOV_LD  ����P}�$PARNUM�  �+?Q�#S[CHy ȕ
�wplq�y��uUPDl�=u���E_CMPa_u����_�'ݥ~%�ER_CHK3��ۣ �G�0�B�RS8A �ȡ_MOp���_���E_RES+_G� ���
��p� "��F�9�j�]�o��� ��ğ���۟����o��@���1��P N�m�r��mP������ ��P̯���`� *�/��f`J�i�n���`�������V 1���ށ�@]s�8��THR_IN�RA �q]مd�M�ASS)� Z=�M�N(�[�MON_QUEUE �������!ބN*�U�n�NkƔȫ�END8��Ώ��EXE������pBE���ϫ�OP�TIO��׋��PR�OGRAM %���%��習��T�ASK_It �O?CFG ��π��ߵ�DATAx����G2�$�6� H�Z�l������������� �2���IWNFOx�혝� ��������������� 	-?Qcu� ������N�Z�� ����pK�_�����z�5G���2�D X,�		x�=��=��@����$a�����0_EDIT ��������WERFL���Ó#RGADJ7 ��AЛ@R$�?�]%0�5&��?�����?�D��A<��z�%�o`�/)(/s#2�'V"	H��l�¾�!?8�Aٴɻt$26*A0/C2 **:L2�??�Q3m=���2�5��+1�9��/�?y= �=�?�?�?�?�?KO�? O5O+O=O�OaOsO�O �O�O#_�O�O___ �_9_K_y_o_�_�_�_ �_�_�_�_goo#oQo GoYo�o}o�o�o�o�o ?�o�o)1�U g������� �	���-�?�m�c�u� ���ُϏ�[�� �E�;�M�ǟq����� ����3�ݟ���%� ��I�[��������� ǯ������	�ߖ� 𰄿����39߿53���ϧ�0�B�o'PREOF �*00�
5%IORITY�:���9!MPDSaP8�'*�"��UT��|34&ODUCT����E��&OG_TG$ ������TOENT 1��� (!AF�_INE��Y�J��!tcpdߌ��!ud{ߴ�!�icm���.��X�Yx#���1)�� Y1�*�0� �S�6�B��f��� ����������!�3���W�>�{���*��x#��)�"�/������BY7/c<��44��(��.A�",  �u�(}���+%��^Ŀf�x�,9!PORT_NUM���0�9!_C?ARTREP% ��aSKSTA�� �4LGSV������#0Un?othing����L�]TEMPG ����T���_a_seiban�,/�</b/M/�/ q/�/�/�/�/�/�/�/ (??L?7?p?[?�?? �?�?�?�?�?O�?6O !OZOEOWO�O{O�O�O �O�O�O�O_2__V_ A_z_e_�_�_�_�_�_��_�_o�VERS�I����M` �disabled�'oSAVE ����	2670H�782J�o�o!`$�o�o���o 	xH��V��.�eK t���J�c|�o����mb_� 1�
���`*�p�!�4��F��W�URGE_�ENBЪ�(���W�Fr�DO���+�W�RГ���WRUP�_DELAY ��,��R_HOT %{���#����R_NORMAL�����W�&�SEM�I6�\���U�QSKKIP���#�xo ��	o��(���Y� G�}�����g�ů��կ �����C�1�g�y� ��Q����������	� Ͽ-��=�c�uχ�M� �ϙ������Ϲ��)���M�_�q����$R�BTIF��0RC_VTMOUE����DCR�Ǿ�� ���5��9C^)C�6�Z@���@�n�6悔���5�O��R������-��>�;�7�� <�	<�S�;�9<���<#*o<���M�Q 7��� y��������/�A��S�e�w������RD�IO_TYPE � ����EFP�OS1 1�ui� xA
-���G2 k�o�*�N�� ��1�Ug N���n�� /�/Q/�u//�/ 4/�/�/j/|/�/?? ;?�/_?�/�??�?�? T?�?x?O�?%O7O�?��?OOjO�O��OS/2 1�ԋZO��O_�O6_�O��3 1��O�O�O,_�_�_|�_L_S4 1�c_�u_�_�_?o*oco�_S5 1��_
ooVo��o�o�ovoS6 1͍o�o�o�oiT�>S7 1�"4�F���"��S8 1Ϸ������~���5�SMASK 1���  �� �NՇXNO���:�<D���MOTE���=�Z�_CFG ��a���A���PL_�RANG]��ߛ�O�WER �%��ΐ��SM_DRY�PRG %%�%�^��ԕTART ��ƞ�UME_�PRO���p�=�_�EXEC_ENB�  ���GSP�DI������Ѣ�TD�B����RMϯ��I�A_OPTION������U�MT_"݀T��_���*�z���9���C�ˀ�����������O�BOT_ISOL�C"�����ֵN�AME %��_���OB_ORD_NUM ?Ƙ���H78�2  ˄h�@�h�$�hʬ�h�>�PC�_TIME�ם�xޏ�S232z�1�����LTEA�CH PENDA1N��v�A�~�]��H@Mainte�nance CoKns˂��ˆ"��DDNo Use ~�E��i�{ߍߟ߱�����NPO#���A��!���CH_LfL��U���	3�~��!UD1:Y�z �R܀VAILI�����U�SR + %������R_INTVAL����������V�_DATA_GR�P 2�%���X�D��P��W���{�f� %��������������� $&8n\� ������� 4"XF|j�� �����//B/ 0/R/x/f/�/�/�/�/ �/�/�/�/?>?,?b? P?�?t?�?�?�?�?�? O�?(OOLO:O\O^O pO�O�O�O�O�O�O_� _"_H_6_l_U��$�SAF_DO_PULS��V���X��QN�PCAN�������SC���(����Gˀq����Px�C�C��˂ p� o0oBoTofoxoo�o��o�o�o�o�o��B���be�!r �dt�:ql�(s�� @���fx��~Ny� �D�t�_ @�T�����~�T D��*� S�e�w���������я �����+�=�O�a��s�����`u2���ǟі��C��¯;�o2���p�����
�t���Di���aC��  � ���Cђax� �Qa�s���������ͯ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ�����������1�2��aZ�l�~� �ߢߴ�������9�u �(�:�L�^�p��� ������2�0�D� �N�	��-�?�Q�c� u��������������� );M_q� ������ %7I[m�� ���D��/!/3/ E/W/i/{/�/�/
��/ �/�/�/??/?A?S? ������r�?�?�?�? �?�?�?O#O5OGOYO gIzO�O�O�O�O�O�O �O
__._@_R_d_v_ �_�_�_�_�_�_�_o@o*o<oNo`o5�艟 9�ko�o�o�o�o�o &8J\n�����pj�o��.2���S�����	123456�78+�h!BO!ܺ�4���`��|�������ď֏ ������o5�G�Y� k�}�������şן� ����1�C�U�f�$� ��������ѯ���� �+�=�O�a�s����� ��h�z�߿���'� 9�K�]�oρϓϥϷ� �������Ͼ�#�5�G� Y�k�}ߏߡ߳����� ������1�C�U�� y������������ 	��-�?�Q�c�u��� ����j������� );M_q��� ������%7 I[m���� ���/!/3/E/W/ {/�/�/�/�/�/�/ �/??/?A?S?e?w?�?�?�?�sm��?�?�q/OO*OF�C�z  Bpqj  W ��h2�bm��} ph
�G�/  	��r2�?�O��O�O�Ook>�_Dlo�<��OB_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o '_�o�o�o�o( :L^p���� ��� ��$�>ISB��1�AiB<S���$SCR_GRP� 1��8�� � � ��SA dE	 ����������1B���SGେۏɏ�:M�4s@��D^@D/^���E��� \ARC� Mate 10�0iD/1450�ҁAM�ҁMD45 678SC
12345��	9��ӅE����KyBד_��SF�߃� S ��Ó��Ӂ�	yJ6��H�Z�l�~�SD�G�H������� ��Əǯ���Ά�oSAگC�֯g�N���v�B�M@Ʋ���ɴ��9A^@ؿ  @S@�f��@��� ?P�Ŭ�HM@)�ۺ��F?@ F�`S�[� ~��jϣώϳ����� ����!ߤ�� �L�7�I�[�m�B�{���� ������	����?�*� c�N��r��_��)������dG�@��0�tSB�@P7H�_D�!�@�p�M@Ȇ�����߃�?��SDAA��������� QƒSA 3E���!ht�U (� ������� �$SF_�EL�_DEFAULT�  ����S@@HOT�STRL��`MI�POWERFL � BEX?�WF�DOM �RV�ENT 1������w L!DUM_EIP.����j!AF_�INEL/SD!�FT�@./d/!����/ �S/�/!�RPC_MAI�N�/�(��/�/�#V�IS�/�)��/H?!7TP;0PU??��d7?�?!
PMON_PROXY�?��e�?�?[2�?�f��?,O!RDM_'SRV-O�gOxOG!R���O�hgO��O!
� M�?�i��O_!RLSY3NC_��8�O\_�!ROS��\�y4K_�_!
CE]0�MTCOM�_�k�_�_!	�RCON�S�_�l�_@o!>�RWASRCGO��m/o�o!�RUS	B�o�n{o�ow/�o ;C�o�o%Jn5�Y�:RVICE_KL ?%�� (%SVC�PRG1����u2��
��p3-�2��p4�U�Z��p5}����p6�����p7͏ҏ�p��$��9�"��t�O J��q�r��q����q G��qo���q��� �q��:��q�b��q� ���q7����`�گ� ������*��؟R� � �z��(����P� ʿ�x������� ȯB�D����r�p� �p����<�������� 	�B�-�f�Qߊߜ߇� �߫��������,�� >�b�M��q����� �������(��L�7� p�[������������ ����6!ZlW �{�������2V�z_DE�V ���MC:��T4���pGRP 2������pbx 	�� 
 ,� ^����/�&// /\/C/�/g/�/�/�/ �/�/�/?�/4??X? j?��?E?�?�?�?�? �?OOOBO)OfOMO _O�O�O�O�O�O�O�O _q?_P__t_[_�_ �_�_�_�_�_o�_(o oLo^oEo�oio�o�o �o�o3_ �o6 ZAS�w��� ����2�D�+�h� O������oy���� ߏ��@�R�9�v�]� ������П����۟� *��N���C���;��� ��̯ޯů��&�8� �\�C�����y����� ڿ��ӿ�g�4�F�-� j�Qώ�uχ��ϫ��� �����B�)�f�x� _ߜ߃�����)��߭� �,��P�7�t��m� �����������(� �L�^�E�����w��� o����� ��6 ZlS�w�������D��d Ԗ�	2{f�`����O%��</�����4!� 4%D/R'</r/`/�/�/ �/�)/�/0)�/?? >?,?N?P?b?�?�/�? �/�?�?�?OO:O(O JO�?�?�O�?pO�O�O �O�O_ _6_xO]_�O &_�_"_�_�_�_�_�_ oP_5ot_�_hoVo�o zo�o�o�o�o(oLo �o@.dR�v� � �$���<� *�`�N��������t� ��p�ޏ��8�&�\� ����L�����Ɵȟ ڟ���4�v�[���$� ��|�����¯į֯� N�3�r���f�T���x� �������:��J�� >�,�b�Pφ�tϪ�� ��Ϛ�ߖ��:�(� ^�L߂��ϩ���r��� �� ����6�$�Z�� ����J��������� ���2�t�Y���"��� z�����������:� 1��
��R�v� ���6�* :<N�r��� �/�&//6/8/ J/�/��/�p/�/�/ �/�/"??2?�/�/? �/X?�?�?�?�?�?�? O`?EO�?OxO
O�O �O�O�O�O�O8O_\O �OP_>_t_b_�_�_�_ �__�_4_�_(ooLo :opo^o�o�o�_�oo �o �o$H6l �o��\~X�� � ��D��k��4� ������������ ^�C����v�d����� ��������6��Z�� N�<�r�`��������� "��2�̯&��J�8� n�\���ԯ������� ~���"��F�4�jϬ� ��пZ��ϲ������� ��B߄�iߨ�2ߜ� ���߮��������\� A��
�t�b���� ����"��������� :�p�^����������� ��� "$6l Z��������� � 2h�� �X����
/� /p�g/�@/�/�/ �/�/�/�/?H/-?l/ �/`?�/p?�?�?�?�? �? ?OD?�?8O&O\O JOlO�O�O�O�?�OO �O_�O4_"_X_F_h_ �_�O�_�O~_�_�_o �_0ooTo�_{o�oDo fo@o�o�o�o�o, noS�o�t�� ����F+�j� ^�L���p�������܏ ��B�̏6�$�Z�H� ~�l����
�۟��� ���2� �V�D�z��� ����j�ԯf��
��� .��R���y���B��� ��п������*�l� Qϐ�τ�rϨϖ��� �����D�)�h���\� J߀�nߤߒ���
��� ���ߴ�"�X�F�|� j������������ 
���T�B�x���� ��h��������� P��w��@�� ����X~O �(�p���� �0/T�H/�X/ ~/l/�/�/�//�/,/ �/ ??D?2?T?z?h? �?�/�??�?�?�?O 
O@O.OPOvO�?�O�? fO�O�O�O�O__<_ ~Oc_u_,_N_(_�_�_ �_�_�_oV_;oz_o no\o~o�o�o�o�o�o .oRo�oF4jX z|���*� ��B�0�f�T�v�� �Ï�������� >�,�b�����ȏR��� N�̟�����:�|� a���*���������ȯ �ܯ�T�9�x��l� Z���~�����Ŀ�,� �P�ڿD�2�h�Vό� zϰ�����Ϡ��Ϝ� 
�@�.�d�R߈��ϯ� ��x����������<� *�`�߇���P��� ���������8�z�_� ��(������������� ��@�f�7v�jX �|����< �0�@fT�x ����/�,/ /</b/P/�/��/� v/�/�/?�/(??8? ^?�/�?�/N?�?�?�? �? O�?$Of?KO]OO 6OO~O�O�O�O�O�O >O#_bO�OV_D_f_h_ z_�_�_�__�_:_�_ .ooRo@obodovo�o �_�oo�o�o* N<^�o�o��o� ����&��J�� q��:���6���ڏȏ ���"�d�I����|� j�������֟ğ��<� !�`��T�B�x�f��� ����ү���8�¯,� �P�>�t�b���گ�� ѿ�������(��L� :�pϲ���ֿ`��ϸ� ������$��Hߊ�o� ��8ߢߐ��ߴ����� �� �b�G���z�h� ��������(�N�� ^���R�@�v�d����� �� ���$�����( N<r`������ ���$J8 n���^��� �/� /F/�m/� 6/�/�/�/�/�/�/? N/3?E?�/?�/f?�? �?�?�?�?&?OJ?L1��$SERV_M�AIL  T5�J@�0HOUTPU}T?H0H�RV 2��6  M@ (�1O�O4D�TOP10 2�>�I d P?�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o����p���5�EYPE`L�NEFZN_CFGw ��5MC�L4oB�GRP 2��%�� ,B �  Ae�L1D;�� Bf��  B�4L3RB21޳FHELL���5��@�O<�ΏK%RSRݏޏ�� )��M�8�q�\����� ��˟���ڟ���7��I�[��  ��+�[�����i��� �L0��ŢơL8q�2�L0d�������HKw 1瞋 ˯ @�J�D�n��������� ߿ڿ���'�"�4�F��o�j�|ώϊ�OMM� 螏�Ϗ�FT?OV_ENB?D�A���OW_REG�_UI��2BIMI_OFWDL����μh�3�WAIT�� ��oE^�Z@��DX�wTIM������VA>@i�3�_UNcIT�����LC�WTRY��4@�MON_ALIA�S ?e���@heOM�_�q��J;� ���������� �2� D�V��z��������� m�����
.��R dv�3���� ��*<N` �����w�/ /&/8/�\/n/�/�/ =/�/�/�/�/�/�/"? 4?F?X?j??�?�?�? �?�?�?�?OO0O�? AOfOxO�O�OGO�O�O �O�O_�O,_>_P_b_ t__�_�_�_�_�_�_ oo(o:o�_^opo�o �o�oQo�o�o�o  �o6HZl~)� ������ �2� D��h�z�������[� ԏ���
��Ǐ@�R� d�v���3�����П� ����*�<�N���r� ��������e�ޯ�� �&�ѯJ�\�n���+� ����ȿڿ쿗��"� 4�F�X��|ώϠϲ� ��o�������0��� T�f�xߊ�5߮����� ���ߡ��,�>�P�b����$SMON_�DEFPROG �&������ &*S?YSTEM*i����<{�R�ECALL ?}��� ( �}7�copy frs�:orderfi�l.dat vi�rt:\tmpb�ack\=>19�2.168.56.1:1968���0�B�T�}.��mdb:*.*�����������_�2x��:1\q�����8 ��,(>Pc�3��a��������d�tpdisc 0�8 ��'9K^��tpconn 0 	��� ]�������./@/R/ e� /��/�/�/�/�� v�/*?<?N?a�/ ?��?�?�?��z/ /&O8OJO]/o/
O�/ �O�O�O�/�/�??"_ 4_F_Y?k?�O�?�_�_ �_�?�?�?�_�_0oBo �_gOo�Oo�o�o�o �Ox_�o�o,>Pc_ �o�_����_�_ |o�o(�:�L�_os� �o����ʏ�o�o� $�6�H�[m����� ��Ɵ��t�� �2� D�W�i����T���¯ U��z����.�@�R� e����������п� ��~���*�<�N�a�s� �ϨϺ���߯r��� �&�8�J�]�o� ߓ� �߶���ۿ�v��"� 4�F�Y�k��Ϡ�� ������|����0�B� ��g����������� ���߀��,>Pc� ���������t� ���(:L_�� ���������x $/6/H/[m/��/��/�/��$SNP�X_ASG 2������!��  0�%y��/?  ?��&�PARAM ���%�! �	*	;P���o4��� OFT_K�B_CFG  ���%�#OPIN_�SIM  �+�j2�?�?�?�3� R�VNORDY_DOO  t5�5B�QSTP_DSB�>j2HO�+SR ���) � &�n:�O��&TOP_ON_ERRO~�FPTN �%��@�C�BRING_PRM�O�#BVCNT_GP� 2��%l1 0x 	DO?_�-_f_Q_�_�'VDPRP 1�C9m0{Q�1m_ �_�_�_�_o4o1oCo Uogoyo�o�o�o�o�o �o�o	-?Qc u������� ��)�;�M�_����� ������ˏݏ��� %�L�I�[�m������ ��ǟٟ���!�3� E�W�i�{�������د կ�����/�A�S� e�w���������ѿ� ����+�=�d�a�s� �ϗϩϻ�������� *�'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ����������1�C� U�|�y����������� ����	B?Qc�u���RPRG_�COUNT�6��B�	ENB�O�M���4�_UPD �1�nKT  
 ��ASe��� �����//+/ =/f/a/s/�/�/�/�/ �/�/�/??>?9?K? ]?�?�?�?�?�?�?�? �?OO#O5O^OYOkO }O�O�O�O�O�O�O�O _6_1_C_U_~_y_�_ �_�_�_�_�_o	oo -oVoQocouo�o�o�o �o�o�o�o.); Mvq����� ����%�N�I�[� m���������ޏُ���_INFO 1Y�/ �� ��R�=�v�a���������*�XEB���C3�B��ƀC!xX�Y?SDEBUG� 0����d��SP_�PASS�B?~�LOG �/�9  ������  ���?UD1:\���_MPC$�/��$��/[�Я /��?SAV �'�����G�_���f�S�VԛTEM_TI_ME 1�'�: 0  �����үr�4�SKM�EM  /�.G�  ��%s����Ͽ��� @��� Q�������"?��׿:A��� p�D�TV���nʟ���� �Ϧϸ���^��E�'V W�������+� =�O�a�s߅ߗߩ߻� ���������{�9� K�]�o������� �������#�5�G�Y��k�}���T1SV�GUNS*�'����ASK_OPTION� /:���_DI�����BC2_GRP 2�/�Q�%���@�C�:��BC?CFG ��s ����`� �������! E0iT�x�� ���/�///?/ e/P/�/t/�/�/�/�/�/?���,!?�/T? f?�/C?�?�?�?�?�? ׮O���0O2O OVO DOzOhO�O�O�O�O�O �O�O_
_@_._d_R_ t_�_�_�_�_�_�_o �_oo*o`oFh10to �o�o�o�oFo�o�o�o "FXj8�| �������0� �T�B�x�f������� ҏ�������>�,� N�P�b�������roԟ ���(���L�:�\� ��p�����ʯ���ܯ � �6�$�F�H�Z��� ~�����ؿƿ���� 2� �V�D�z�hϞό� �ϰ��������ҟ4� F�d�v߈�߬ߚ߼� ������*���N�<� r�`�������� ����8�&�\�J�l� ���������������� "XF|2ߔ ����f� B0fx�X�� ����///P/ >/t/b/�/�/�/�/�/ �/�/??:?(?^?L? n?p?�?�?�?�?��? O$O6OHO�?lOZO|O �O�O�O�O�O�O_�O 2_ _V_D_f_h_z_�_ �_�_�_�_�_o
o,o Ro@ovodo�o�o�o�o �o�o�o<�?T f���&��� ��&�8�J��n�\� ��������Əȏڏ� ��4�"�X�F�|�j��� ����֟ğ����� .�0�B�x�f���R�� Ư������,��<��b�P���p���A���*SYSTEM*���V9.0055� ��1/31/2�017 A v�  ��K�TB�CSG_GRP_�T   \ $ENABLE��$APPRC_�SCL   �
$OPEN�C�LOSE�S_M�INF2'�ACC|��PARAM�� ���MC_M�AX_TRQ��$d�_MGNk�C��AVw�STAL�w�BRKw�NOL�Dw�SHORTMO_LIM�ʧ�h�9J����PL1��6����3��4��5��6
��7��8k�q���?� $D�E��E��T��b�PA�TH^�w�m�w�_R�ATIOk�s�T� �2 	$CN�T�A�����m�I�NX�_UCA�~��CAT_UM���YC_ID 	����_E����6�������PAYLO�A��J2L_UP�R_ANG6�LW�A�?�3�O�x�R_F�2LSHRTv�L�OD���}��Ӌ���ACRL_S�ؽ����+�k�HVA�$yHx���FLEX���J2� �P�B_F��$^��_FTM��&���$RESERaV�>�;�� ����� :$���LEN.�z�;�DE|���;�Yғؔ���SLOW_AXI^��$F1��I���2��1������MO�VE_TIM��_?INERTI��
��	$DTORQCUEX�3��#I��ACEMN��%E�%Ep	V��d�A8�R�TCV��@Rt����
��T@�RJ���	�M��,��J_�MOD����� �dRy�2��P�pE���\�X���AW�gQJKh@��K��VK�;VK�JJ0����JJ�JJ�AA6��AA�AA%�3AA �t�N1�N �d�#��E_NUv�� g�CFG�� � $GR�OUPc�SK��B�_CON�C��B�_REQUIRE����BU��UPD�ATT�EL�}  �%� $kTJ��� JE��gCTR��
TN �F�&�'HAND_kVB��OP�7 $oF2x�3��m�COMP_SW��ѣ��R�� '$$Ma�e�R�Î8����<� �5�¼6A_�.�h�D�<q�A��A���A��A���0��D���D��D��P��GR�ǂAST�ǂA���AN��DY���x� �4�5A���s��s��2�B��R����P ����� �)�2�;��#� �0i�\�� 7�U6��QAS�YM��
�TС�p�мݎ���_SH�" �������TU8����%�7�J>���P�pcfi\o�_VI83�h|6þ`V_UNI���d�{�JU�bU�b ���d���d v���� ������su��� �@��HR_T��a	N2�q���DI���O�t�p�#
)  �2I�QAz��� �q �S�s � g� ��p  � f1MEe���pr�QT�pPT&`r a�>���~$�5`C�^��R�T4`! $�DUMMY1�o$PS_ RF��֤�$����FL�A� YP_��F�?$GLB_T�0�u�΅>���g�; 1�qc X��'�STf�� SBRv�M2�1_VT$SV_ERa�O(`�,�SCL��Ap O�r��pGL�`EW�� 4 $H�$Y�2Z�2Ww��x�Bb3A��Ҥ�W�U]�� oN��)`w$GI0}$]�� d�W���� qLh���'b}$F'b�E��NEAR_ N��F�\ TANC���<1JOG���� �e�$JOI�NT�& ��MSE]T�  ��E畄� S��˕� ���  Ue?��� LOCK_F�O��m1�pBGLV�3GL��TEST�_XM�j�EMP�=�Ϣ悖�$1UC�\���2� ��B����i0������CE| Ó� $K�AR�M�sTPD�RA`�3�*�VEC�~�D�.�IU���!C{HE��TOOL���i�V��REK�IS�3;���6���AC)HP���v�O��F����29���I�� � @$RAIL__BOXE�� oROBOƤ?��?HOWWAR���<����ROLM��ŀq!��¡!Ӱ��J�O{_F� ! �����K�6��pRN�OBo�6���?�C��Y�OUR������Q�"�!��$PIPǦN]�Ӳ�� ���V�@�CORDEAD����u��p� O�p  D ̀OBA�#�������p̀��'`�!SYS���ADR�!�p>�TC}H�0  ,oSEN�r#�A��_���d�z!��AC�pV�WVA� �� 9�]��uPRE�V_RTA$E�DIT��VSHW�R�!�&��]q���`D(�.Q��6Q$HEAD8amp�КHa��KEq�|�C�PSPD�JMP��L�uV�Ra �tQ���\�IРS�"�C20NEr��!�'T'ICK���QM�QjR�:�HN�� @p�W�~%�_GP��ʶ$�STY^ү�L�O�<2:���� t 
��Gj�%�$�Ѳ�=��S�!$�aJp-����p��9P�P��SQU-���<���aTERCB�gR��TS�$  ����']�'-`�>p1OC�6�bPIZ��������PR�������S��PU�a��_DYO�c�XSN�K�v�AXI��/���UR� p�"찕�"�]1�� _`�4�ET5P(��ЦU��F�W��A�A�Q��ĳ���!5�g�RE4lu��9��:��6�	 �2��7��9��9� G�G�'F"TI�F�R&��4C�E o2oDoVd�!SS}CЀ  h� cDS��4���SP�p&"%AT@�2����c⅂ADDRESzs�B��SHIF�#^�_2CH� ѹI�t!�TU�I�1 6�CUSSTOV��V��I�rA UҸ�6!��P
Ϫ�
�V������! 	\��������,��J�2CSC��Y�*��2��1�TXSCRE�E��"�p�TICNAO���T4����866"vP# TI�/� ��4�.���63��4��RRO�@�3а
��1�6�UE?�$# ��PMѧ�SP�4��RSM����UNEaX_�vA�pS_���+F�SA.IIG�S6Cx��B�4 2#O0UErT%�r?�nF��WGMT3pL�a��O@��BBL�_��Wo���& �����BO���BLE�f"�C밚"�DRIG�H�CBRDA�\!C�KGRo�UTEX�$ UQWIDTH�����Ʊ��Jq 7�UI>�EY6 ��' dh��Ѐ���Ӱ=��BACK�ᡂ4�UE�!�FO���W�LAB�?(!�I<����$UR��P��_P'�H�1 ( 8wq�_��t"�R(�Rq�����������R�QOm!��)��L��PU�@7cR���L�UM7cV ERVH��D�_PP�fT*�j GE�R�a `�M)�LP�e_E\���)�g��h!�h����i5�k6�k7�k8 �bZ�6����4�������SJ�)^QU{SR]�+ <��b'�U���#��FO� .��PRIrm��%qވpTRIPϱm��UN�p�t,�� ��p������]P�3 �-� -�RSp��G  �T/��u!�rOSF��vR9 �2�so���.f�x�����$���U�a��/$�6�pDC�b���sOFFŠ���0��L�O�� G1.9�����/9�GU.�P���׃��sQSUB��H��@'SRT��1����;���OR��'�RA�U� (�T=�Z��V�C� Ҕ2� ɲ��$���y�8��`C��{�DRIV��@_V���������D4tMY_UBY3t�����$��19��l0��	����P_aS�����BM�A�$b�DEY_�E�X�@�3����_MUb.�X�An� @USA 8��p[�k0w�xp� �2�x�GgPACINr�!�RG�𦥽���`��A���SCp�RE�R�j!o��`���S�3{ � TARGÐ!P72���a�R�S�A4nP0`TQ�	o����REz�SW��_IA��� o���OIq�\!An v��E$pU��෱� \Pa�HK
��5����y��s�̦0��EA��ɷWO�R�Pv����MRC]V�A6 ��`O��M�PC83	����REF�G(���� e�s`cM�Xp�^���^�-ˀ�Ƶ�_RCʻ���0S!pf�ϓ���Lma��D7 �@��gPTU0 epԕw��OU�����惓 S2��2 $U00��r�45#�^��K SULb�5fc`CO�0 `6`� ]��Ӥ0���Ѫ�a��@q��i�L���$��՘a��@q�s�?�8�| +5#k� �5#CACH��LO R�&�<�a�A�KQC ��C_LIMIg#F�Rj�Tl���$H�O�P�*�COM	M��BO�@��ب �a��VP��/ ��	_����Z����k����WA{�MP�FA�Ik�G��;�AD<?�p�IMRE�_���GP@V�� k�A�SYNBUFk�V�RTD������&SOMLo D_|���WA��P�ETUO�X�Q�����ECCU�V�EM٠%�k�VI�RC?����B��_DELA����p�p��AG��Rc�XYZM@5Cc�W3�qsQ� T��P��qs��D9�"�QLASAP�
�� Gl� :�rX�S�a�7�N�_�LEXEE�;�3W�ka5!���FLPIW���F�I����F���P�:#�<_p�
���8t@s���@ORD�|qȎP��##�� =*_0Z`T�r�B�1OJP6b �SFE �3�>  a0s���c�U�R�⟱SM�u?ȬrV�R J� f���"�5@�r��qL�IN��@�WN�X�S屎 A��2��K�&SHd`HOLk���XVR�t�B��@T_OVR~k �ZABC��C��"q-1  ��Zހ�tD�rDB�GLV��Lϒ�R��ZMPCF�E��0�t2ޑLN�~ ��
m1d��F� Ђ`��ɰ4CM�CM��C��CAR�T_Y1��P_2` �$Jw3q4D ��}2�2�7`�5`��sUX|5UXEu��6|�5�4�5�1�1��9�1�6����Z�%G`*�$W�AuYV D�p H�R1RM�{qy�HET��$��PU'�Q��@>�I � �3��� PEAKf���K�_SHI�B��'R�V F^`G½B� C �@r2g1|�����A20ұ�I S��DXTRWACE�PVw�	A�SPHER'aJ� ,e�THjO|I��$TBCSG� �2 @�Q������ � ` �_�_�_�_�_�_ �_�_.ooRodkwR~S��\d ���a?�Q	 HCB�do�iC  B `�R�o�h�o�kB��o$p��o�jdf  AXp?�w{qW �{������@�@�:nT�g�z�E� W��������
����3�	V3.�00�R	md4�5�	*U�M��0��1�� ��m���  ��֟�wQJ2{c�]6����n  �U�QY ����E�ş�p��p�����	 _�ȯ���ׯ���4� �D�j�U���y����� ֿ�������0��T� ?�x�cϜχϬ��Ͻπ������>�P�X� 7�j�|�&ߜ��߬��� ��	���-��Q�c�u� ��B��������� ��U%�7��Q��=�c� Q���u����������� ����)M;q_ ������� 7%GI[� ��������/ /�M/;/]/�/q/�/ �/�/�/�/??%?�/ I?7?m?[?}?�?�?�? �?�?�?�?!OOEO3O iOWOyO�O�O�O�O�O �O_�O__/_e_S_ �_w_�_�_�_�_�_o �_+ooOo=oso�o// �o�o5/ko�o�o 9'Io]��� u�����5�G� Y�k�%���}������� �׏���1��U�C� e���y�����ӟ���� ��	��Q�?�u�c� ��������ͯ��� �o�oA�S���+�q��� ����ݿ˿��%�7� I�[���mϏϑϣ� ���������3�!�W� E�{�iߋߍߟ����� ������A�/�Q�w� e����������� ���=�+�a�O���s� ����e���������' K9[]o�� �����#G 5k}��[�� ���//C/1/g/ U/w/y/�/�/�/�/�/ 	?�/-??=?c?Q?�? u?�?�?�?�?�?�?�? )OOMO_O��wO�O3O aO�O�O�O�O__7_ %_G_m__�_O_�_�_ �_�_�_o!o3oEo�_ ioWo�o{o�o�o�o�o �o�o/SAc ew������ ��)�O�=�s�a��� ������ˏ�O	�� -�׏]�K���o����� ��۟ɟ���#�5�� Y�G�}�k�����ůׯ ������1��U�C� y�g�������ӿ���� ��	�?�-�O�Q�c� �χϽϫ�������� �;�)�_�M߃ߕ�?� �߿�i������%�� I�7�m�[�}����� ��������!��E�/��  e�i� �i�}�i��$TBJ�OP_GRP 2�1�� _ ?�i�	��ڜ����9� � ���V�� ��������i� @e��	? �CB  ��C����5GU	i��C 2BH  �A�/��D!�,��bB* qh�$�7C�� A���c�d���i�A �EG +��a	���D/�D<Ky/�//#/�/�/��	??�/ �/T?f?%?o?a	�?�? �?�?�?�?�?O)OO !OOO�O[OO�O�O�OP�O�O_g�i�1Q��E	V3.00���md45���*[P��d�i_tW �G/� G7�� G?h GG8� GO Gd�� Gz  G��� G�| G�:� G�� G��� G�t G�2� G�� Gݮ� G�l G�*� G�� HS��RF� F@� F+� FK � Fj` F�� F�Q � G�X �R�Q^� G�v G�ĨS��4 G�� G��� G�\ G�� =L��=#K�
]Ae�Js�Yokbi�oo�o���ESTPAR�P�]����HR�`AB_LE 1	��C`%i��h�g ��di�g�hn i�h�p�g	�h
�h�h�ei��h�h�hDa�c'RDI�o���o !3EWu�tO��{@����+��bS��� �z����"�4� F�X�j�|�������ğ ֟�����0�B��� Āȏ���g��l�~��� ��N`r���x�b~i�NUM  1����	 q� �C`D`�b_CFG �
R���@��IMEBF_TT�ap�����`��VERBc�������R 1��k 8f_i�dd�� P���  � ��%�7�I�[�m�� �ϣϵ���������� !�3�|�W�i߲ߍߟ���������A�����ƜMD3�E��� 8k�}��V_I���INT�����T1�#�5� B��O�a����_TC������$0�P����9�RQ��RԴ_L���@˵�`MI_CHAN��� ˵ nDBGL�VL��˵�aq E�THERAD ?U�e� ��`������hq ROUmT��!P�!#�ASNMASK��˳�255.�GS}��GS�`O�OLOFS_DI��P�%�	ORQC?TRL ޻7��o-T/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?s</�?��?�?�cPE_DE�TAI��PGL�_CONFIG �R�b���/�cell/$CID$/grp1�?@4OFOXOjO|O2��
 �O�O�O�O�O_�O%_ 7_I_[_m___�_�_ �_�_�_�_�_�_3oEo Woio{o�oo�o�o�o �o�o�o/ASe w�*��������}�O�a�s����������?я��� ���*�<�N�`�� ��������̟ޟm�� �&�8�J�\�n����� ����ȯگ�{��"� 4�F�X�j��������� Ŀֿ������0�B� T�f�x�ϜϮ����� ���υ��,�>�P�b� t߆�ߪ߼������� ��(�:�L�^�p�� ��������� ���@�User� View "I}�}1234567890C�U�g�y���`����. C����)�26���+=Oa����0�3��������	h*��4 �cu�������5R/)/;/M/ _/q/��/��6/�/ �/�/??%?�/F?��7�/?�?�?�?�?�?8?�?��8n?3OEOWO�iO{O�O�?�O�B �lCamera4�*O�O__)_;_M_+�E�Ow_�_�^ A��_�_�_�_�_o)  �F���O_oqo�o �o�o�o`_�o�oLo�%7I[m�O� �F�	����� %��oI�[�m������ ��Ǐُ돒�wQ�� 7�I�[�m����8��� ǟٟ$����!�3�E� W����w+k🥯��ɯ ۯ�����#�5�G��� k�}�������ſl��E �)Z��!�3�E�W�i� ��ϟϱ��������� ��/�ֿ�wm9��{� �ߟ߱�����|���� �h�A�S�e�w��� Bߤw!I2������� /�A���e�w�������������������9 ��HZl~��I� ������ 2DPVhz	J	�E0  �����/�3/ E/W/�{/�/�/�/�/ �/|��@�Ky/.?@? R?d?v?�?//�?�?�? ?�?OO*O<ONO�/ �EBk�?�O�O�O�O�O �O�?_*_<_�O`_r_ �_�_�_�_aO��{Q_ oo*o<oNo`o_�o �o�o�_�o�o�o &�_�U��or�� ���so���_ 8�J�\�n�����9�U ��)�ޏ����&�8� �\�n���ˏ����ȟ ڟ������U򻕟J� \�n�������K�ȯگ �7��"�4�F�X�j��  ����� ��Ͽ����)�;�<M�_�   o�w� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w�����������c��  
�(  }荰( 	 �� ;)_M�q ������%:��� ̹�j |������� /�Y6/H/Z/�~/ �/�/�/�/�//�/?  ?g/D?V?h?z?�?�? �/�?�?�?-?
OO.O @OROdO�?�?�O�O�O O�O�O__*_<_�O `_r_�_�O�_�_�_�_ �_oI_&o8oJo�_no �o�o�o�o�oo!o�o "ioFXj|� ��o���/�� 0�B�T�f�������� �ҏ�����,�s� ��b�t���͏����Ο ����K�(�:�L��� p���������ʯ��  ��Y�6�H�Z�l�~� ��ׯ�ƿؿ�1��  �2�D�V�hϯ��Ϟ� ����������
��.� u�R�d�v߽Ϛ߬߾��������;�@  �#�5�G��� ���0frh:\�tpgl\rob�ots\am10�0id\arc_�mate_��_1450.xml� ������������0�B�T�E���Y�~��� ������������  2D[�Uz��� ����
.@ WQv����� ��//*/</SM/ r/�/�/�/�/�/�/�/ ??&?8?O/I?n?�? �?�?�?�?�?�?�?O "O4OK?EOjO|O�O�O �O�O�O�O�O__0_ GOA_f_x_�_�_�_�_ �_�_�_oo,o>n`��� �k�<�< i�?� >k�o>oyo�o�o�o�o �o�o�o5-O} c���������1�?��$TPG�L_OUTPUT� I�I� a`i�~����� ��Ə؏���� �2� D�V�h�z��������ԟ���
��i�a`��6�2345678901A�S�e�w��� ����?�>�ʯܯ� � �$���(�Z�l�~�����:�}��Կ���
� ϴ�ƿR�d�vψϚ� ��DϺ�������*� ��8�`�r߄ߖߨ�@� R�������&�8��� F�n�����N��� �����"�4�����j� |���������\����� 0B��Px� ���Xj� ,>P�^��� ��f�//(/:/L/�A�}\a�/�/�/�/�/�/�-@co?#?�ij ( 	  &�X?F?|?j?�?�?�? �?�?�?�?OOBO0O fOTO�OxO�O�O�O�O �O_�O,__<_>_P_�_t_�_4��_`xf�_ �_�]�_o*ooNo`o .��_�o�o=o�o�o�o �o!o%W�oC ��y��3�� ��A�S�-�w���� q���яk������ =�����s�������� ������a�'�9�ӟ %�o�I�[�������� ��ٯ#�5��Y�k� ɯS�����M�׿�ÿ ��}��U�g�ϋ� ��wω���1�C�	�� ��'�Q�+�=߇ߙ��� ����i߻�����;� M��5���o���� �����_���7�I��� m��Y������%��� ����3i{ ����K�����/�R�$TPOFF_LIM �P|��Q���JN_SVN  ��$`P_MOoN �Ub���2�%JST�RTCHK �U`/hVTCOMPATu�d�VWVAR r�"(y �� :/Y�J_�DEFPROG %�%Q/�/f�_DISPLAY�U�j"INST_�MSK  �, ��*INUSER���$LCK�,�+QUICKMEN"?ެ$SCREA0��U "tpsc@�$�!\0a9`r0_v9�ST�`RACE_CFG ��"$Y	C$
?���8HNL 2y*�P�1)+ O"O'O 9OKO]OoO�O�O�J�5ITEM 2K� �%$1234567890�O�E  =<�O_*_2S  !8_@[L �O�_C#�O�_
_�_ �_@_�_d_v_?o�_Zo �_jo�oooo*oDo No�oroDV�oz �o�o|&��
� n����:���� ����"�ʏF�X�!�|� <���`�r�֏����L� ՟0��T� �&�8��� D���ҟ�^����گ �P��t������4� ί�������(�:�� ^�ς�B�Tϸ�j�ܿ ����6���ߎ� ~ϐϢϼ���@��ϖ� ����2���V�h�z��� ��J�p���ߎ�
�� .�� �d�$�6���B� ������������� N� r���M��h�� x���8J\ ��,Rd��� ���F//| $/��{/��/��/��/0/�/T/f//?�4S��2�?4:�  �B4: �1�?�)
 �?�?�?�?c:�UD1:\�<���F1R_GRP �1�K� 	 @� :OLK6OlO ZO�O~O�O�N��@�O��J�A�?_�O7_"U?�  R_d[N_�_r_ �_�_�_�_�_�_�_&o oJo8ono\o�o�o�o��o	5�o�oD3S�CB 2P; =_:L^p�����:<UTOR?IAL P;�?��?7V_CONFIG  P=�1�?��?t�$�OUTPU�T !P9e�����ď֏���� �0�B�T�f�x����� b���ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϷ�������  ��$�6�H�Z�l�~� �ߢ߳����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������� �&8J\n �������� /"/4/F/X/j/|/�/ �/�/N�`����/?? &?8?J?\?n?�?�?�? �?�?��?�?O"O4O FOXOjO|O�O�O�O�O �?�O�O__0_B_T_ f_x_�_�_�_�_�_�O �_oo,o>oPoboto �o�o�o�o�o�_�o (:L^p�� ����o� ��$� 6�H�Z�l�~������� Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ������Ͻ(����������6��/Z� l�~ߐߢߴ������� ��� �2��V�h�z� ������������
� �.�@�Q�d�v����� ����������* <M�`r���� ���&8I \n������ ��/"/4/F/Wj/ |/�/�/�/�/�/�/�/ ??0?B?S/f?x?�? �?�?�?�?�?�?OO ,O>OO?bOtO�O�O�O �O�O�O�O__(_:_ L_]Op_�_�_�_�_�_ �_�_ oo$o6oHoY_ lo~o�o�o�o�o�o�o��o 2DS{�$�TX_SCREE�N 1"�;���}�S� ������B� �1�C�U�g�y���� ���ӏ���	���� ?���c�u��������� 4��X���)�;�M� _�֟蟕�����˯ݯ �f����7�I�[�m� ������,�ٿ��� �!�3Ϫ���i�{ύ� �ϱ���:���^����/�A�S�e��ω��$�UALRM_MS�G ?sy��p ��Vj��������"� �F�9�K�i�o����������SEV � �����E�CFG $su�}q  Ve@��  AJ�   B�Vd
 ��]csu }����������������1?&�GRPw 2%0� 0Vf�	 g����I_�BBL_NOTE� &0�T���l]bxp_a�<�DEFPROx��Z�� (%�� _`�*N9r ]��������/�FKEYDA�TA 1'sys �p ?�Vf  =x/�/� g/�/�/�%,(/�/Vd�/?8ANCEL(?S??�w?^8EXT ST�EP�?�?�?�?�5ORE INFO�? �?O*OONO5OrO�O kO�O�O�O�O�O_�O�&_8_ ��/�frh/gui/�whitehome.png9_w_�_�_�_�_��_�_�_o�o,o>o�UFRH/�FCGTP/wz?cancelb_|o �o�o�o�o�_�o�o�0BMo_cnextko������o � ��$�6�H�S]cinfoq������ ��Џ����*�<� N�ݏr���������̟ ޟm���&�8�J�\� 럀�������ȯگi� ���"�4�F�X�j��� ������Ŀֿ�w�� �0�B�T�f�=_uϜ� �������������,� >�P�b�t�ߘߪ߼� �����߁��(�:�L� ^�p��������� �� ���$�6�H�Z�l� ~�������������� ��2DVhz� �����
� @Rdv��) ����//�</ N/`/r/�/�/%/�/�/ �/�/??&?�/J?\?�n?�?�?�??[�;}�JP����?@�?�=�? O2OF,_ cO_�OnO�O�O�O�O �O__�O;_"___q_ X_�_|_�_�_�_�_�_ o�_7oIo0omoTo�o �o���o�o�o�o! 0?EWi{��� @�����/�� S�e�w�������<�я �����+�=�̏a� s���������J�ߟ� ��'�9�ȟ]�o��� ������ɯX����� #�5�G�֯k�}����� ��ſT������1� C�U��yϋϝϯ��� ��b���	��-�?�Q� ��u߇ߙ߽߫����� �o��)�;�M�_�f� �����������~� �%�7�I�[�m���� ����������z�! 3EWi{
�� �����/A Sew���� ��/�+/=/O/a/ s/�//�/�/�/�/�/ ?�/'?9?K?]?o?�? �?"?�?�?�?�?�?O �?5OGOYOkO}O�OO �O�O�O�O�O__���![������J_\_n]F_�_�_|V,�o�_�o�_�_o -ooQo8ouo�ono�o �o�o�o�o�o); "_F�j��� ������7�I�[� m�����O��Ǐُ� ���!���E�W�i�{� ����.�ß՟���� ���A�S�e�w����� ��<�ѯ�����+� ��O�a�s�������8� Ϳ߿���'�9�ȿ ]�oρϓϥϷ�F��� �����#�5���Y�k� }ߏߡ߳���T����� ��1�C���g�y�� �����P�����	�� -�?�Q�(�u������� ��������); M_������� �l%7I[ ������� z/!/3/E/W/i/� �/�/�/�/�/�/v/? ?/?A?S?e?w??�? �?�?�?�?�?�?O+O =OOOaOsOO�O�O�O �O�O�O_�O'_9_K_ ]_o_�__�_�_�_�_ �_�_�_#o5oGoYokoh}o�of��k�f�����o�o�m�o �f,�C� gN������ ����?�Q�8�u� \�������Ϗ���ڏ �)��M�4�q���b� ����˟ݟ��o%� 7�I�[�m���� ��� ǯٯ������3�E� W�i�{������ÿտ ����Ϭ�A�S�e� wωϛ�*Ͽ������� �ߨ�=�O�a�s߅� �ߩ�8��������� '��K�]�o���� 4����������#�5� ��Y�k�}�������B� ������1��U gy������� �	-?Fcu �����^�/ /)/;/M/�q/�/�/ �/�/�/Z/�/??%? 7?I?[?�/?�?�?�? �?�?h?�?O!O3OEO WO�?{O�O�O�O�O�O �OvO__/_A_S_e_ �O�_�_�_�_�_�_r_ oo+o=oOoaosoo �o�o�o�o�o�o�o '9K]o�o��@������ ���� ����*�<�N�&�p���\�, n���f�׏������ 1��U�g�N���r��� �����̟	���?� &�c�J����������� ����)�;�M�_� q��������˿ݿ� ϐ�%�7�I�[�m�� ϣϵ��������ό� !�3�E�W�i�{ߍ�� ������������/� A�S�e�w����� ����������=�O� a�s�����&������� ����9K]o ���4���� #�GYk}� �0����// 1/�U/g/y/�/�/�/ ��/�/�/	??-??? �/c?u?�?�?�?�?L? �?�?OO)O;O�?_O qO�O�O�O�O�OZO�O __%_7_I_�Om__ �_�_�_�_V_�_�_o !o3oEoWo�_{o�o�o �o�o�odo�o/ AS�ow���� ��r��+�=�O� a����������͏ߏ n���'�9�K�]�o��F q��F ��������������̖,ޯ#�֯G�.� k�}�d�����ůׯ�� ����1��U�<�y� ��r�����ӿ����	� �-��Q�c�B/�ϙ� �Ͻ���������)� ;�M�_�q� ߕߧ߹� ������~��%�7�I� [�m��ߑ������� �����!�3�E�W�i� {�
������������� ��/ASew� ������ +=Oas�� ����//�9/ K/]/o/�/�/"/�/�/ �/�/�/?�/5?G?Y? k?}?�?�?x��?�?�? �?OO&?COUOgOyO �O�O�O>O�O�O�O	_ _-_�OQ_c_u_�_�_ �_:_�_�_�_oo)o ;o�__oqo�o�o�o�o Ho�o�o%7�o [m����V ���!�3�E��i� {�������ÏR���� ��/�A�S��w��� ������џ`����� +�=�O�ޟs�������л�ͯ߯�0��>�0���
�� .��P�b�<�,Nϓ� FϷ���ۿ�Կ��� 5�G�.�k�RϏϡψ� �Ϭ���������C� *�g�y�`ߝ߄����� �?��	��-�?�Q�`� u���������p� ��)�;�M�_���� ����������l� %7I[m���� ����z!3 EWi����� ����///A/S/ e/w//�/�/�/�/�/ �/�/?+?=?O?a?s? �??�?�?�?�?�?O �?'O9OKO]OoO�OO �O�O�O�O�O�O_�� 5_G_Y_k_}_�_�O�_ �_�_�_�_oo�_Co Uogoyo�o�o,o�o�o �o�o	�o?Qc u���:��� ��)��M�_�q��� ����6�ˏݏ��� %�7�Ə[�m������ ��D�ٟ����!�3� W�i�{�������ï R������/�A�Я e�w���������N�㿀����+�=�O�&P�Q��&P���zόϞ�v����Ϭ�,��߶�'��K�]� D߁�hߥ߷ߞ����� �����5��Y�k�R� ��v���������� ��1�C�"_g�y����� ����п����	- ?Q��u���� �^�);M �q������ l//%/7/I/[/� /�/�/�/�/�/h/�/ ?!?3?E?W?i?�/�? �?�?�?�?�?v?OO /OAOSOeO�?�O�O�O �O�O�O�O�O_+_=_ O_a_s__�_�_�_�_ �_�_�_o'o9oKo]o oo�oX��o�o�o�o�o �oo#5GYk} ������� �1�C�U�g�y���� ����ӏ���	���� ?�Q�c�u�����(��� ϟ������;�M� _�q�������6�˯ݯ ���%���I�[�m� �����2�ǿٿ��� �!�3�¿W�i�{ύ� �ϱ�@��������� /߾�S�e�w߉ߛ߭ߴ�ߖ`����`����������0�B��,.�s�&��� ~����������'� �K�2�o���h����� ����������#
G Y@}d���o� ��1@�Ug y����P�� 	//-/?/�c/u/�/ �/�/�/L/�/�/?? )?;?M?�/q?�?�?�? �?�?Z?�?OO%O7O IO�?mOO�O�O�O�O �OhO�O_!_3_E_W_ �O{_�_�_�_�_�_d_ �_oo/oAoSoeo�_ �o�o�o�o�o�oro +=Oa�o�� �������'� 9�K�]�o�v������ ɏۏ�����#�5�G� Y�k�}������şן ������1�C�U�g� y��������ӯ��� 	���-�?�Q�c�u��� �����Ͽ���� ��;�M�_�qσϕ�$� ���������ߢ�7� I�[�m�ߑߣ�2��� �������!��E�W� i�{���.������������/��$UI�_INUSER � ���P���  �0�4�_MENHI�ST 1(P�  (_���(/SOFT�PART/GEN�LINK?cur�rent=men�upage,153,1o�����s�)����631��pew�� �'-?95T�����8�k}��������� / /$/�H/Z/l/~/�/ �/1/�/�/�/�/? ? �/1?V?h?z?�?�?�?���D1��D?�?�?O O)O;O>?_OqO�O�O �O�OHO�O�O__%_ 7_�O�Om__�_�_�_ �_V_�_�_o!o3oEo �_io{o�o�o�o�oRo do�o/AS�o w������?�? ��+�=�O�a�d�� ������͏ߏn��� '�9�K�]�o������� ��ɟ۟�|��#�5� G�Y�k���������ů ׯ������1�C�U� g�y��������ӿ� ����-�?�Q�c�u� �ϊ��Ͻ�������� ��)�;�M�_�q߃ߕ� $߹���������� 7�I�[�m��� �� ���������!���E� W�i�{�����.����� ������Se w�������� +��as� ���J��// '/9/�]/o/�/�/�/ �/F/X/�/�/?#?5? G?�/k?}?�?�?�?�? T?�?�?OO1OCO.���$UI_PA�NEDATA 1�*���yA�  	�}�  frh/cg�tp/flexd�ev.stm?_�width=0&�_height=�10�@�@ice=�TP&_line�s=15&_columns=4�@�font=24&�_page=wh�ole�@UO1) � rim�O!_   �@8_J_\_n_�_�_�O �_�_�_�_�_o"o	o Fo-ojo|oco�o�o�op�o�o�o1� @r/_4FXj| ��o�%_���� �0�B��f�M���q� �������ˏ����>�%�b�t�[���| ��{C�۟����#� 5���Y��}������� ůׯ>������1�� U�g�N���r�����ӿ �̿	��-�?ϲ�ğ uχϙϫϽ���"��� f��)�;�M�_�q߃� �ϧߎ��߲������ %��I�[�B��f�� �����L�^��!�3� E�W�i��������� ��������A( ew^����� ��+O6s ���������/ /h9/��]/o/�/�/ �/�//�/�/�/?�/ 5?G?.?k?R?�?v?�? �?�?�?�?OO�� UOgOyO�O�O�OO�O F/�O	__-_?_Q_c_ �O�_n_�_�_�_�_�_ o�_)o;o"o_oFo�o �o|o�o,O>O�o %7I�om�O� �����d!�� E�W�>�{�b������� Տ������/��S��o�o}�d�������ӟ���)����u� H�Z�l�~�����	�Ư ���ѯ� ��D�+� h�z�a�����¿Կ������x�c�k�$UI�_POSTYPE�  �e� 	 �[�*��QUICKMEN  9�H�^�,��RESTORE �1+�e � �뿑r�����ϑrm �)�;� M�_�q�ߕߧ߹��� �߀���%�7�I��� V�h�z��ߵ������� ���!�3�E�W�i�{� ��������������� ��Sew�� >�����+ =Oas(�� ��//'/9/� ]/o/�/�/�/H/�/�/ �/�/?�?0?B?�/ }?�?�?�?�?h?�?�? OO1OCO�?gOyO�Ox�O�Oi�SCREy��?~�u1�sc��u2�D3��D4�D5�D6�D7r�D8�A�CTAT5��� ���e"�US#ER�@�O�BT�@�CSks�C�T4�T5�T�6�T7�T8�Q*�N�DO_CFG a,9�t�s�*�PD-Q�gY�No�ne *�^P_I�NFO 1-�e`��0%�O,o�x o[o>oo�oto�o�o �o�o�o!EW�:{b��QOFFS�ET 09�a �PC��XO���� /�&�8�e�\�n��r� ����ȏ�����+�"��4�F����ϒ�����
���ڟ�xUFRAM/E  PD�V�Q�RTOL_ABRqT���s�ENB�~�GRP 11�����Cz  A� u�s��Qs��������� ͯ߯��x�U?��Q~.�MSK  B��a.�N��%	i��%b���k�VCMRv[�27�{#��R@	�Pfr1:� SC130EFG2 *ݿ�PD���Y��T&��5R@�Q�?��@�p���N�� ɟ5�?� IH`�rϟ�ı����8�-�A�RB����RB B��� �RA#ի�Dߋ�h�7� ��w߰ߛ��߿���
� a���@�+�=�v�)ߚ���ISIONT�MOU�B��U����R8S�߸S� j� _FR:\��\�P�A\�� �� wMC�LOG�   UD1��EX5�RA' ?B@ ��x�I��r���I����PC �� n6  ����IFu�%���`��Z�  =�C��PD	 J�*�TRAIN_���nǐ  dPp	�栲9�}(c�� W������� .2@Rdv�Z��_\�RE��:b��ʲ��LEXE��;ܪ{�Q1-e��VM/PHAS/P�U�S�Ж�RTD_F�ILTER 2<.�{ Ԓ��,�{/ �/�/�/�/�/�/�/? ?��i/N?`?r?�?�?��?�?�?�?�?��SH�IFT�1=�{
 <��q�JODU)O OO�O_OqO�O�O�O�O �O�O_<__%_r_I_�[_�__	LIV�E/SNAPes?vsfliv.�_W��� �pU�P�Rmenu�_�_�_ Woio@b	E��>IO�VEMO��?�� ���$WAITDI�NEND��+��dO ?�"��g���oS�iwTIM@���<|G�o^}�o�{az/xazN�hRELE%!�@��d�����a_AC�T�P�K�E�� �@d�ko���E�RD�IS�PA��`V_A�XSR�p2Ab������Vp_IR  �j 	��)� ;�M�_�q��������� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��������XVR�a�B��$ZABCvp1C� ,N rf�2ϵ�ZIP��D�e����������MPCF_G 1Eٍ0J��=���S�FىX�`# �c�߆�<90 ��߻�S�|��ߠ�?�}������S��$��z�8���� �����������
�4��M���G��JÛ�Y�LINDK!Hً� Є� ,(  *��������������� ��);M ��p���{�� � U6��l S�w�����Y�s2Iه]� �)� #/3,���\/G/�/��h/�/���!A�c��SPHERE 2Ju��*?z�/<? #?`?��/�?�?$�? k?Q?O�?&OO?\O nO�?�?�OO�O�O�O��OEO"_4_F_M�ZZ/� ǘf