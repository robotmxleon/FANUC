��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A   �����
�WVAMP_�T   �$X1  $kX2AY@  /�FC5  �$2ENBA $�DT T_R�2 d ENA�BLEDnSCH�D_NUMA  �/ CFG5�� $GROU�P�$z ACCE�L@�G$MA?X_FREQ�2 �L�DWEL�D�EBUG�PRE;WSOUT��PULSEAS�HIFt 7TYP�4$USE_A�EF} 4$GD=O�  f0� r?�NpW�EAVE_TSK� �V�_GP��SUPPORT�_CFnCNVT_DONE p �}k}GRP #2r�� _� ��$� TIME1�o$2'EXT�� (1#&(MODE�_SW�CO3 S�WIT �/ PH�AX6  4 �� ECC$�T�ERMNnPE�AKno!AL � \ � �!I֑$�!N_VSTAR�#!r"ؾ�"�%�CY�CL42 
ISST/ � Tv"b �$CUR_RE�L_� �!TW�PR5 � 
�$CEN� _RI�3RADIU��XIz ] Z�IMUTi!$E�LEVATION�g5� N�CONTINUOe2q �MoEXAC=PE����1�6  H|~ �UENCYA��ITUD4�2RgIGHC�2LEB�L_ANG1 ��OTF_� ?	�  $3A�bET��n3C!$ORGjH�FBKjH��P���C��DLDW�HR�E�_�3�B�C��D��B�C�@�D�A�CCHG�G	Q�F	Q�F	Q�FINC�G=Q�F=Q�F`=Q�F�AVCPYC� _T�\#�Y~P#�@�SY��H)@�U�PD"0n�$$�CLASS  ����Q��8 �P��PVERS�1�W�  ��~�QIRTUAL�_��Q0 2�X�{ �   ?��@�  HaDae�T Woio{o�o�o`)dNw 2 3k Hf���uHe@O߀Hi�oNc)a� � e�� E`��H��$���
��2  �z����=�����4s ����jpYq��w�r��Dq��x at��ujp`��i.�5t8q�q2�b�t���
�<q`����� @q����̏ҏ���Sb�)a�  23k
=TDaSI�8�� �����Cph�?m�'R ����l�D��� ��Ca��l����k���� �2�D�V�h�z��l�FIGURE 8��o�v�Hal� f��������M�(� H��󈯎�����Ŀֿ~�TCIR1��Pd�}�0�~�h�0z�D�Z�l���0�v� ��~����� ��$ߪjN� Hp��4q�Ȓ���@��ʖD�M` g����������	���-�?�Q�c�u�`�� �q� �5)�ᐟN`���ᬟ ����˟���M�_�q�������������k�Triangle��z�h߾�M�� Ɵ�ύ�����0�/ L� &��g�n�� �	//-/?/Q/c/u/ �}DVhz��/�/ ��9?K?]?o?�?�?�?�?�?����� O �h��O2ODOVOhOzO �O�O�O�O�O�O�O
_ _.[�?._O"O�_�_ �_�_�_�_�_oo&o�8oJo\ono�mSCH�EXTENB  �=��ctSTAT�E 2�k �|o�o�o �gWPR 7�6�L}D��-�_OTF 	8��@)0�q�q����v)��uAȫs�u@�  <#�
�?�����mu_GP 2w| ���d� v����я㏡+