��   F��A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A #  �����#�AMON_D�O_T   �$PORT_�TYPE  �@NUMJ/SG�NL7 L�$MIN_RAN}GI$MAXr�NOo ALxp V��~ �COUNT>J��AWE08 �� $AWn0ENBJ $�|G1LY_TIV�$WRN_ALM�STP�
�E��C�.�WT�C�
J�AFT_�CHGxAVRG�_INT��{SgAVE�YP1?ER_REG�Tw$WA� SIG�� OP��V/OLTS�����AMP�&AEx �#E_VL� �&D'>% I*f$� _�ANL�  �p 
$US0 S�_CMD � PRIORITY�"�UPPER� $�LOW�$�#$FgDBK�"�RAv ~�!SQ_AVG�#n�#SD_� CE� 8� ��$ �� � �LIN�!$ARC_ENABL�!|� 0DETEC�!~< ELD_SP�$?PD_UNI��!N92DIS�"�ID sIM�#�� � v1WFt2 ����CF�" � �$PS_MAN�UF �2O�DEL�5PROC�ESN0�0WFEE�W0ESC�2�2_F�I#1�1�1�7T _A�O�"�2I�6D�7D�C1�6L �"{2 ι CNV� 7 ?  $EQ�zlxODOU�θ�?@TBd  �$?C 2 �kEDD   �, � MM�!�$D� ��!?2 $F� �B�kBE?@7	JBSE�L10_NOJDA�TA_s@�@ VkBWPpG
{M
�F;WP7 L@�L�
 �WIR_wCLP4 L@�ASBU8  H �$4��Rx�4�YPREF� <�U�_ECU�� � JB~ �S _  $BPEEP�f#}!SCH7 � �!��`��1e#dPK*jFwREQ.gULSwbSP�0fg2y�!hyb*g�FZ b06 �ZCoVG}�h p dD�e�e�`�	�a���dBVB�aZERqOy}uSLO]R�`NT�!P�cO	U\�93�L FORMA�0NAra�0J3	� D�cQWUX�WEIOEX7O4 �A�Wfx�ccpS_91IN�p� :1�U�p� FcAUG"t0LO�0�qP�!�G��R<�yADp;�STIC�@��pROBOT�A{DY�rERRO�SE��`S��p�!�TR��$S�CHD�OG_�@%��0_AOCTIV���I��C�01�2�q�O�TF7 � $
��P��x�nfpNCi0�c;� f0�*d;�*g0�7f;� 7i0�Fd;�Fg~�Td���TfUP�@�B�#PC�R7�� WS#TK��� =�Hr Ւ Ɓ%��00��2�X���0A~�3KIPTHE91�S;������PIKEf���0��0WWV�2t�E_�HO;0�0��PHKp-1���� RMT����SPTL�0p�3$Hz��SW��pd�$BBg1_ONL4�$B�2pf�bgF�WF�1e2_R`��zE"�!� _W;6~�AND1OFF��.�!ND2g�3g�R��S� �A� 9CEPM~� | $�0 �@g��e��*f��7b���Ff�TfADAP�T� G�CSENS��c��!ݒ��8 � 0?,2���"� �$�1b�!c�7cc�Fa |�Tac�^��'y��&l�T�&�!4�&5�&6�"p8�W�@�2 HOU�!��o � �SE �0�g4�Q�T<��6 �'��46�q56�0� %$CURR7�(��"HEATzP e@�!燰"j���i�p.��GAP�#Ti�XP�Y0��EHP��@��pDYS�@�!GP�0S�!�$���$GO� RI���AM�#/"�#�M��jAN3O�BE	FB ;�LHV1[5j�@�43;1 `H�V�PA�H�r���3��F1�� ��DPOSR 7� � 	� RSB �$��0G�m�b�O�J�X��O��DU�IW�"AXQl�2C,1LB�"D����?3|!E��8  4�@P֋q]ִSGʦ�~�;A8�~8  $ $�@��CL�$��s	�P|��8 $ ;o2 � �"�ql��q��� 	PK�P��
��*�� �q�Ba��b�@4�5�6:2K�`3�����FW�q��B��ALAR ���2��2����t�
�3�Q_R}���
�.44�F�+�P	W,���_@ĸ�Ӕ ]�������Qbw0m��t���QDI�c��j��~pus�R�SIyZ���BOAR��D�1]E7�]�\ �h"0h"��ķ�_$VEND��I��DEVIC��0D\����MAJ��V�#�IN�(�$�uI"�vM1A��pFI�0�B�W��RE�� p $��X�� ⡡��MF̀OR_R��C��^1D4TO_��O5_�R�pRS�Q'�OS܇9�qEUP� #N��S�0�`�=�� �6��6��9PUcRG��RKtSTF!R�p&���A��.E �.E�AED��P-��	M%�fMT�����eEM7��Q�5���Z$�2 2�9�P駇��K�p�Q�ADJ�T��NEX�T��r_LE�c��P��X��M����aA�B�_�#IV���H�q��2�eFL������P ��U���0�8� ��T�WT[�CY�� ���  ��	`��`( �bTOT�AL_�Q�c���VI�p�WWARo��U��A*�PY&1b�uKG���'" A}�#�N�p  ��SwCFG�1z��LOO�B:��P�Q��S!@���GLO�B�P�⣠� ��NO-T��$0QI4�*��AVh�Y��$���������e��W_S+HFL�W�X�fkr�I�$�q �e�RY�	��оP��%�ʀLI�MS`�i�@�c7�UI�F�e�APCOU�PL�R @ ��p�q��� �qU�R�`N��<�MM�Ym �u0�u�  �����USTOk� ?   x�0 ��qp` 
,�SEsMGg��1! ,��cMG�Ag���NOzP�R ����wa�"� ,/���Ȣ=6 Ƞ��3T� )�RT����p�=����AHE R�A�������'"݈ {�������@���Q� L��)BD ��2C���x7B<�i3_FIL@��W��BUG_3SM ���ñF_F����hq�, _4N SV@Ђ�TC�P��=Ҕ�DIO�������.af�TM�C��PA�P�q��qw�x��q�_DYNV�2Wԣ����KEYV�GQׂ���F��?�/B�{�_uC��R�TOU��p���Б��CAL�Q�0�`� TIp1�P_Fy�RT���@��A?2���$$CLA�SS  ��e��� ��� ��-�SB����  ���IR�TU�����AWA�OY1�� 
���$�
�K���n�29�f�[�[���g�
�?������� g����������� (�:�L�^�pςϑ�l�EXEu�`������� ��Ͽ�*�<�N�`�r���ߖߨߺߕ�r@S Rw���:����#� 5�G�Y�k�}��������������n�N�LG 2x� �����?��<1�6�`�	�e��� p`����{`� 2:�)��Genera�l Purpos�e�MIG �(Volts, �0)��� ����
�AWMGENL.�VRA*EG�LMG19��g� `��������'���� ���������~�CNV 2	x�{�[���.�� 4aPz Uh�����/ /�=/O/./s/�/\ �/�/b/�/�/�/?'? ?K?]?<?�?�?r?�? ��E�/�?O�?2ODO #OhOzOYO�O�O�O�O �O�O
__�?@_R_�O v_�_g_�_�_�_�_�_ �_o�_(oNo�?ro-_ �o�o3o�o�o�o �o8J)nM_� {o������ � F�%�j�|�[������� ֏�go���0�B�!� f�E�W���{���ҟ�� ����,�>��b�t� �������ί௿�� ���:�L�+�p���� O���ʿU�� �߿$� 6��Z�l�KϐϢρ� ���ϯ���ߵ�2�D� #�h�z�Yߞ�}ߏ�������
��NVWP� 2|	i\>�T� 
��b�t���USTOM 2|l  ��������h�	hd"���D�EFSCH R|�Q�<�b�@�Default Schg���n����� ������K" 4�Xj��������
)�FBKL�OG1 @��T�῀  Ugy��12=O�����5LG_CN�T  ����)�I�OEX 2������A ��C�]$@������!�
�Weld Spe�e%��IPM  d$�/�/�/�/??�(?:?��OTF 2��A?�?�?�?x�?�?C8=������@����?K)�PC�R 2��pI�B	H�?��BDCN<D7�������?�ffAAZ �A"��OFM"@����/�O@uO"@����9��OELG��k%*_��F�02345678901JRG��A%4_y_�_�_HIȩ_|7]�OOSRAM2���IB�$�_oCRGSEL R<��Q� 	Pro?cess 1oRSf2�_oj3i�o4i�o5�-mlXSJ���o7��kn8i�'l"@��� c�_);Es-B� ��W�%Vol�tage��qs�fc%Dw|!@]�y�h��a�Wire f�  s�$	� hc%[& t/�oDS�l*�<�N� `�r���������̏ޏ�����&�]+zvd"�����  �#��E�Z"!��a��^/>�� ��V���a��aɒCurr�ent�Amp �=���l�eu���Q� c�u���������ϯ� ���)�;�M��W�� �a�����ឱ	q��)q ��Iq��R�͹ϧg�a �aA��b-���-�	q-��)q-�ZU!��\e��	q?�����Z �%������ϻ�����8�PDRuS R\zH���jq��C�U�g� ����gߩ߻�u߇ߙ� ��������]�o�)� ;�M�������� #������k�}�7�I� [�����������1 C��I��Wi ������?Q /����� �//)/;/M+�U/ g){/�/�/M/�/?cS2
�S^=R��b�S2�UPYp^=�=��o?�33H1>>E0=L��>I0hU!�"�#�$�1Lt9�g�q�#?�v�#>�8�8CWIR/E 2&M<�?�?�h�>�3�>��G(=�J*�ES?CFG �G�A ��Y��OOˎE7])C�OUPL�0=k
0�vkB`�D�^�L �[�OZW�O�G_�OP_�G_Y\�HNB  ���Ec&FUSTOM  =k
8ƙy�O�&EEMGOFF �!=kS��)BP�CR "�_�@	���zqC{sUūMJo@�\zt�f_oeo��
Cl �q¨1