��   v1�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����UI_CONF�IG_T  � E$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY6]5�ODE�
6CWFOCA �7C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"�%�!BA�!j ��!�BG�#�!hINS�R$IO}7P}M�X_PKT?$IHELP� {ME�#BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�<ST]Yf2$Iv!_Gv!k FKE�E ��8C�&USTO}M0 t @;AR$@PIDDbB�ChD*PAG� ?�^DEVICEބISCREuEF���}GN�@$F7LAG�@�KB��1  h 	$P�WD_ACCES � =EFB�S:1~�%)$LABE� O$Tz j�@��32R�	�CUSR�VI 1  < �`'R*'R�(QPRI�m� t1�P�TRIP�"m�$�$CLA�@ �����Q��R��R̜P\ SI��W  �׸QIRTs1�_�P'2 �L17�L1A��R	_ ,��?���b�P$c ca��� , ��  Ao��
 ���'/SOFT�Pb@/GEN�1?�CURRENT=|>�A,18,1lo��o�o�o�o �o�o,95,2�o?QcNu �(5�` w�����)q9�G�Y�k�}��� �s�oˏݏ������E,381�oN�`� r�����Q������ӟ ���	���-�?�Q�c� u��������ϯ�� ���)�;�M�_�q������aTPT�X��&���˿`� s����$/s�oftpart/�genlink?�help=/md�/tpmenu.dg��2�D�V�h�!� �Ϟϰ�������u�
� �.�@�R�d���uߚ� �߾������߃��*�`<�N�`�r�����Q�[f=fc��($ ��������������Qa:�<o��F���A���zc��\a���^�����  ���	���������8�8�]�:�W` � ��� ���SQB 1�XR_ \��_�� REG �VED��FXw�holemod.�html	sing}l}doub��trip�?brows�t� Y��CUg�y��C-gyd/ev.s�l/� 1,	t0/�/ ��/�/�/m/�/�/p�/�/?8?� �P P?b?t?�?�?�?�?�?�?�?�6 @L?!O3O OWOiO{OJF;	3?-? �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_�oo3oEo Woio{o�o�o�o�o�o �o�o/ASe wE?������ �0�B�T�OOx���Y� k���ҏ�O�O��� '�9�b�]�o������� ��ɟ�����:�5� G�og�a�������ů ׯ�����1�C�U� g�y���������ӿ� � �2�D�V�h�zό� �ϰϫ����ϵ���� .����ݿv�q߃ߕ� �߹��������%� N�I�[�m����q� ��������!�3�E� W�i�{����������� ����/��j| ������� �0B#x�A� S�9����// '/9/b/]/o/�/�/�/ �/�/�/�/�/��?? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�OY�O�O�O�O _ _2_D_V_h_c�_��_m__�_�_�Z�$�UI_TOPME?NU 1�Pa�R 
�da�A)*de�fault�O�M�*level0{ *�K	 Ho�60�o/o�o�btp�io[23]-8?tpst[1�h�o��o�oko}o(=h5�8E01_l.p�ng</6mencu5^yUp�q13^z�r]z}t4�{l)q����
��.�@�R� �B�{�������ÏՏ~d�prim=�q�page,1422,1܏�'�9�K� ]�h���������ɟ۟�j���class,5��+�=�O�a�l���13h������¯ԯ�m���53��"�4�F�X�j�m���8�����ɿۿ� l��#�5�G�Y�kϖI`a.o��Rm��+q0������fty�m�o��amf[0�o��	>�c[164�gf�59�h+q�ߣ�yx2��}�ҙz��w]{ ��s����n���� ����������"�4� ��X�j�|�������A���2����/A ���w����N `�� $6H��	�1\������M���ainedi��//)/;/M/H��config=single&��wintp��X/�/ �/�/�/�Ja���/? Se?%��E?W?i?|? �?�?�?�?1?�?�?O O/OAOSOeOwO��O �O�O�O�O__M�>_ P_b_t_�_�_'_�_�_ �_�_oo�_(oLo^o po�o�o�o5o�o�o�o  $�oHZl~ ��1�����  �2��V�h�z����� ��?�ԏ���
��.��N��d����������O��5�s�̟�'�ٗuݤ��� �����@3��ڂ�����̩6ٯu7�F�X�1�C�U� g�y�ď������ӿ� �����-�?�Q�c�u���f"\1k���� ����	��-�?�Q�c� u߇�߽߫������� ��Z�M�_�q����$�6�6��������0��d$�74$�U� g�y������,C���5�	TPTX[20196��4��246�������18"4(F��0�25��10��i���tvԡ�H���0�1����C:l$treeOviewy#�3C�&dual=o�81,26,4$ �����////A/ S/e/��/�/�/�/�/d�/&�;x�53� �E�O?a?s?~/�?�? �?�?�?�?�?O'O9O@KO]OoO�/?:�1%?ª2���O�O�O �y6�O.�edit� �O�OT_f_x_'�w5� 1_CS�_�_�_o��o 4o�<o�Uo!{o�o �o�o�o�o�ogo /ASew��� �����"�4�F� Oj�|�������ďS� �����0�B�яT� x���������ҟa��� ��,�>�P�ߟt��� ������ί]���� (�:�L�^������� ��ʿܿk� ��$�6� H�Z�	oo��?o�� �������� �1�C� U���aߋߝ߰����� ����	��@�R�d�v� ������������� �*���N�`�r����� ��7�������& 8��\n���� E���"4� Xj|����S ��//0/B/�f/ x/�/�/�/�/oρ��/ ��?���=?O?a?s? �?�?�?�?)?�?�?O O(O9OKO]OoO1�O �O�O�O�O __]/6_ H_Z_l_~_�__�_�_ �_�_�_o�_2oDoVo hozo�o�o-o�o�o�o �o
�o@Rdv ��)����� �*��N�`�r����� ��7�̏ޏ����&� �/�/\�?���?�O�� ��ǟٟ����!��� -�W�i�{�������ï կ�O��0�B�T�f� ��x�������ҿ��� ���,�>�P�b�t�� �Ϫϼ������ρ�� (�:�L�^�p߂�ߦ� �������� ��$�6� H�Z�l�~������ ���������2�D�V��h�z���:�H�*d?efault��j��*level8��M��	�� �tpst[1]�	KyPtpi�o[23R6Hu�P����me�nu7_l.pn5g��13�	�5
��41u6�
�w���� ���//+/=/O/ �s/�/�/�/�/�/�/~n"prim=��page,74,1�/?-???Q?c?n"��&class,13h?�?�?�?�?�?u?�25�?"O4OFOXOjOm#|<O�O�O�O0�O�O�/218?)_@;_M___q_|O�26x_��_�_�_�_�_��$�UI_USERV?IEW 1J�J��R 
��EDIT,�Weld DAT�A s�doub�lej���_�medit1eo�o�oh�o�okj�&95P �o,>�o�ot����p�0cSTATUS,POS@ftripMo_oqo��,�>�P�b��Yy2�m�����ÏՏx�33 _��1�C��P�y� t������˟ݟ�� ��%�7�I�[�m���� ����ǯٯ�����
� |�E�W�i�{���0��� ÿտ���Ϯ�/�A� S�e�w�"��ϖϨ�� ������+���O�a� s߅ߗ�:߻������� �ϸ�"�4��X�� ������l������ #�5���Y�k�}����� L������D�1 CU��y���� �v�	-?�� L^p����� ��/)/;/M/_// �/�/�/�/�/v�/�/ �/n/ ?I?[?m??�? 4?�?�?�?�?�?�?!O 3OEOWOiO?vO�O�O O�O�O�O__�OA_ S_e_w_�_�_>_�_�_ �_�_o�R