��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����DRYRUN_�T  4 �$'ENB  �$NUM_POkRTA ESU@�$STATE }P TCOL_���PMPMCmGR�P_MASKZE�� OTIONNLOG_INFON�iAVcFLTR�_EMPTYd ?$PROD__ L ��ESTOP_D�SBLAPOW_�RECOVAOP�R�SAW_� G� %$INI�T	RESUME�_TYPENDIST_DIFFA $ORN41� 8d =R ��&J�_  4 u$(F3IDX��_ICI  �MIX_BG-yy
_NAMc �MODc_US�d�IFY_TIv� �MKR-�  $LI�Nc   "_SIZ��� �. �X $USE_FLC 3!�8:&iF*SIMA7#�QC#QBn'SCAmN�AX�+IN�*}I��_COUNr�RO( ��!_TM�R_VA�g#h>�ia �'` �����1�+WA-R�$�H�!�#�N3CH�PEX�$O�!PR�'Io�q6�$$CLAS�S  ���Ԕ1��5��5�0VE�RS��7�  �ץ1IRTU� �?�0'/ �5_5��������0F�0�1E��%�19O��5OnO������5I2�; !�O�O�O�O__'_ 9_K_]_o_�_�_�_�_`�_�_�O+ W?�8�0 ��j�0�*o<oNi�� � 2��9  4%�_�o��AA�o�o �o�o�o%7[��@�AM�=��p�����dcs�y@jc$"+ uk"K�0��1U�A`�XA�1 �0$N��������Џ� ���*�<�N�`��� FAu�A������ʟ ܟ� ��$�6�H�Z�0l�~��4L�a�C�7 2ulu�ۯ ����#�5�G�Y�k� }�������t�ͯ��� 
��.�@�R�d�vψ� �ϬϾ�ɿ������ *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx �������� ,>Pbt�� ������/(/ :/L/^/p/�/�/�/�/ �/�/�/rv