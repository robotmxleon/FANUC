��   K�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_���$$C�LASS  ������D��D�VERSION�  ���/IRTUA�L-9LOOR� G��DD<x$p?�������k,  1 <D
wX������ Z)/;/Z�/o/�/@�/a/�/�/�/_ �/��/	?';�$MNU�>A�  <���d?/\<t5s?z';�3C��ד? y?�?�?�?O�?O3O aO)cO�OwO�O�O�O �O�O_�O_E_�;5�NUM  ���x�S0tUTOOLC?o\ 
Y8]��2}?��;�.�TP/3��4�R��P�Po¨�m�2��V IO[_oCOoAo'o9o [o]ooo�o�o3_�o�o �o�o#EsY {������X�V y�Wy