��  U��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A0  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ����AIO_CN�V� l� RA�C�LO�MOD�_TYP@FIR��HAL�>#INw_OU�FAC� �gINTERCEmPfBI�IZ@�!LRM_REC�O"  � AL]M�"ENB���&sON�!� MDG/� 0 $DEBUG1A�"d�$�3AO� ."��!_�IF� P �$ENABL@�C#� P dC#U5K��!MA�B �"�
f� OG�f d PCOUPLE, �  $�!PP=_D0CES0�!e8Y1�!"PC> Q�� � $SO{FT�T_IDq2�TOTAL_EQf� $�0�0NO�2�U SPI_IND�E]�5Xq2SCREEN_NAM� {e2SIGN�0�e?w;�0PK_F�I0	$TH{KY#GPANE�4� � DUMMYE1dJD�!UE4RA�!RG1R� � $TIT1 d ��� �Dd�D� �DTi@�D5�F6�F7�F8�F9�G0�G�GPA �E�GhA�E�G1�G ��F�G1�G2�B!S�BN_CF�!	 8� !J� ; 
2~L A_CMNT�$FLAGS]��CHE"� � E�LLSETUP �
� $HOM�E_ PR<0%��SMACRO�RR'EPR�XD0D+�0��R{�T UTO�B U�0� 9DEVIC&�CTI�0�� �0�13�`B�Se#VA�L�#ISP_UN9I�U`_DODf7{iFR_F�0K%D1�3��1c�C_W�Aqda�jOFF_�U0N�DEL�hL�F0EaA�a7b??a�`$C?��PA#E1�C#sATB�d�� W_PL�0CHn/ <� PU�P"�B
2ds�`QgdswDUT�PHAgp�SF��WEL�DH2/0 =pLc7w7atAING�0�$�r�1�@D2�4%$AS_LIN;t�E�w�t_��2UC�C_AS
BFAI�L�DSB"�FA�L0�AB�0�NRDY��P�z$��YN�Wq<��`DE 6r��`���+�����tSTK��+�;s7�;sNO�p��[�̈́r��U* Ȁ%�9 � � � ��q`�G�C�G�+�U�S_FT�vpF�ǂ�G�SSF��PAU�S���ON7xǓHkOU�ŕMI�0�0ƔSEC�2�ryi �rHEK0�v8vGGAP�+�	�I� Ν GTH���D_I���T= �l�� ���`�s9!̅����9!G�UN1���q���#�MO� �cE �� [M�c����R�EV�B7���!X�I� �R  �� OD�P-�	�dPM���%�;�/�"8�� F��q�P1X�0DfT �p E RD_E�%�Iq$FSSB��&$CHKB�pEFdeAG� �p�  "H
�Ա� Vt:5��8�3 a_EDu � � C2��q�S�`�vl �d$O�P�0�2�a<�_OyK��Y�TP_C� �<�d�vU �PLAC��^}��p� xaCOMM� �rD|ƒ��0��`�KO]B�IGA�LLOW� (tK�w�0VAR��d!�1}#BL�0S �� ,K|aԚPS�`�0M_O]=՗_�CCG�`N�!� �� ��_ID_��� �0�� B.��1S� ~�CCBD	D�!��I�����@�Ҍ84_ CCWp�` OcOL
��P'�MM
�zn�CHs$MEAdP��d`T�P�!��TR1Q�a�CN���FS3��ir�!/0_�F��( D�!��
`C�FfT X0GR�V0��MCqNFLI���0UJ�����!� SWIl�&"D�N�P�d��pM�� � �0EED��!��wPo��`�PJedV
�&$�p�1�``�P��ELBOF� �=��=�p/0���3P�� ������G� �A0WARNM�`ju��wP��8�𼠤 COR-��8`FLTRjuTR�AT Tlp� $7ACC�rTB� ��>r$ORI�.&ƣ�RT�P�pg=m��CHG@I��"3�T{�1�I �r�  3 K���� ����"�Q���HQD���a�2
BJ{P�C��3�4�5��6�7�8�96�COfS_rt�����3�V�OLL�EC��"MULTI�b
2��A
1���O�0T_�R ; 4� STY2�R
���).��p�P0m� |A06Kb�Ib$���Pc����UTO=�cE�EXT!Y�
B!�Q? 2 
l��a0��Rub����  �"�� �Q����qc�o~#A!|��1Y�M
��P8$  lTR>�� " Lq��/���P��`AX$J�OB׍��b� 5IGx# d��?%? 78��3�p%��Lq�CO_MOR��$� t��FN�
CNG&AF�TBA���6 �JC��9��D@r��1CUR.KPa`/E^ ,�P��%��?��t�taoA��XbJ��_R��|rC�LJ�r�H�LJ�DA���I�����2G����RfT&� ��byG���HANC6$LG��iqda��N��*�YaCᇁ�0|rf�R
'L��mTX���nS3DBWnSRA�SnSAZ`�X��$  ' gFCT��e�_F��IPn�e�M
P�QIkOh������1��e� ���Cg���A���cMPa� ��HK�&AEUp�p�Q�2 9 ��'  ]PI>��CSXC��ZqG( xs��s��T�R��CcPN����MG��IGH"��aWI=DR�$VT�P�Ŗ9�EF�PA cI��XP,aQ�1u�CWUST��U��)R"GTIT����%nA[IO����P_�9L���* \q���OR��$!�q���-��OeP��jЅpIp �Q�u�J8�
��0��� @ DBPXWO�RK��+[ $S�K0���v"BT)PT}Rw� , �l@AAb��s�R0�ؠD��A:0_C����=�+`FH�PL�q��R�A�"D��#�D��r����ȑBJ���9��� &] DB�Q��-�r~q�PR��ΰ
�D8ct��. �E�\S�a���LӉ/����( ��0�R�P�j� 1%�b��rA�E���� 2D��b�W��RE���3�HPC�  7.$L��/$Ӄ������INE׶�q_9D����ROS��E�0"2q��f0�p��P�AZ�tAsbETURYN����MRQ2UA@v�CRŐEWMwp^��SIGN�A&r�lPA��W�`0{$Pf1$P�P&�2j���q������DQ��f����|��׶GO_AW;0ऱ�vp��qam�gDCS'���CYx	42O�1�8�8���2��2�N�@��C�tDۣDEVIѐ 5 P $SRBֳ��I�P.�i�I_BY�q���yT�A9�HNDG��6�������b�DSBLr3ͳ�7��Le7 H x�� ��TOFB���FEБg')��ۣ�f8��DO�a�� MC9�"�`�sr�(�
�H�PWp�v"ݡ�SLA4���9IINP!Ѐ� ж�ۡ�_:D *�SP Np�#�lƍ�1��W�I1��J��E�q87r�qW��NTV#r��V ��SKI�STE^��b��pڥ�a�J_�Sjb_>���S�AF�k���_SV>BEXCLU��p�o�D�pLX ��YpH��%q��I_V9`�bPPLYj��������_ML��>L�VRFY_D��M�IO�`  P�%`țb�Oe��LS(�|b��4}����	��P�u���Y�AU NFzf�����)���cD�4Ͱ� �S��r�AF� CP�XЁ��&`� ;�j��pTA#��� s ���SGN��<��<@3�P��c_�t��a���qd��rt��`UN>�����<@rD�p]�T`����%`�����9�p�pI>�= @b��F��\t6@OTS� ���|������孁|p[EMr�NIC>2�K�GM A��iDA=Y�sLOAD����D��5��W�EFV pXI�?j����~cO� 7�5�_RT;RQU�@ D�����0Q�p �EԠ��� ?K�%>`|� ���AMP*Pp��A�"'; DB'L��VDUS�U���CABU�B`�N�S9@ID�1WR�$�Q!`V[�V_8#� ; �DI@J$C� /$VS�SE�T�BDC�A� `���|�DB�AE_��;VE�P�0SW!�!�@x�3�� �@�`�OH�@P�P <IRwqDBB �p�=�!U����t"BAS��o'~P�Pn%[�d� B	� ���oRQDW]%MS� ��%AXC'�;LI�FEC���� ��	2N@1EB5��3EBCd@�/Ź�Cq`ʡN0�4q�6��OVՐ%6sHEh�DBSUP�1��	2D�_�4j�H1�_!C�5š�7Z�:W��:qa�7�S��"BX�Z�PʁEAY2HC"��T�pސ�NM��� ��CT�dgD `L��@HE�VXCSIZ?6k0��[��Nh�UFFI�0���C��������6ܭ�zrMSWJEE �8��KEYIMAG�TM���S�A5���F��
q�BOCVI9E �qF 	�P�LQ�_��?� 	���&`KDG� ��ST��!>R|�FT���FT� FT� FPEMA�ILb �aA���FAULSHR�*��;pCOU_��q|pT���U�I< $d�S_�S#�ITճBUFkG�kG@�jpJ`p�0B�Tk�C�p�Rws�PSAV(e �R�+Bd�$ Cg�p��AP/d_ň�$̰_�Pec �iOT�����P@����jA�gAX��sq:p�P��\c_G�3ЁYN_e!�pJ�0Df�W�r�d"M�O_0T��F�����E2���^ЈqK��ey&^�5q9�)�4��qL���nq�S&�cC_ܐ��K씐pu�t��R�A�u�XnqgDSP�FnrPC�{IM5c�s�q�nq��U�w{0�0��PIP�R�nsN!D  �tT!H��"ûr� Tߑ�s�HSDI�vABSC_�9@`�V��x�v���c~����NV��G ��~�*@�v�PF!�`ad�s0p�a��SC��\��sMER��nqF�BCMP��mpET��⌐M�BFU�0D�U�P?�M�B
�CD�yH��`�SlpR_N)O�ዑN� %�i�Xcg��PSf�C?�%v�C���a��d��`U OH����c  d�������}�锍� �9疗疢疮A*�7�8�9�0T��1��1
�1�U1$�11�1>�1K��1X�2f�2���2�
�2�2$�21�2�>�2K�2X�3f�3R�3��
�3�3$�U31�3>�3K�3X�94f�BAEXT�TP <sK�p<6p��p2ǋ��QFDR^�QT�PV���b	2p�v�	2REMr�F��0BOVM�sz��A��TROV�ɳDT3`��MX��I�N��Q0�ʶIND����
	�i��`$DG�a{#��4P5�9D���RIV"�=2�0BGEAR�qIO�K��;N0p}ة��(���@�0<Z_MsCM@	1 �F|0;UR"�R ,t� a�? P0�?\��!?��EG���*Qa��e�S j�!P�a�RIM��P�SETUP2_� T � �STD 6���<����I�C�[���QBACrU T([ �RTt)Nz%��+p�IFIQ!+p���А��PT{b?���FLUI1TV g� Y�PUR�! �W2�r<qv��P�� �I��$�S��?5x#�JQpCOw`�c�VRT� x$S�HO���SASS�Y��a?58����AZ�W�RFU��15q�2fu��*@�X �|�NAV�`��3���*@�R=1���VISIJД�SC����E�c�\�AV���O��B%E�X$PO��I�\ �FMR}2b�Y o� X�}p�bpNt�{ߍߠ�߶ơP���_f�DG�_��B��M4�|Y�k�DGCLFR%oDGDYLD��B7�5!6.�04��MR��3SZ�P�	 T��FS�`2T[ P�!��bs�`$EX_���1�`Ā\2j�3�5��G��J9\��
���PWe}O�&DEBUG��L"��GRR�spU惷BKU�O1�� 0PO� ;)' ���' Mb�LOO��ci!SM� E7bA� ���� _E �] �@Y���T�ERM�%^�%�QO�RIBq� _�&��S�M_OpL� `�*A��)a�%��UPRb�� -���](�#0^��G:0�ELTO{Q$U�SE��NFIc1�G2��!���$4_$wUFR��$j�0A1}0=�� OT�7���TAX�p��3NST�CpPATM�d@�2P'THJ�;�E4P_bD�H2ARTP`R5�P8Pa{RG1REL�:�aSHFT?�H1�1�8E_N�R�8��& � 	$�'H@a�q�B��N�bSHI@�U��= JaAYLO��a �a���Y�1��~�J�ERVA�3H� �7Cp�2�����E�����RC�~�ASYM.q~�H1WJ[7��AE��1Y�>�U2T@Cp�a�5�Q=��5P�X�@��bFORCpMK&a�GRz!:c��'"�`&�0w0�aG_�H9Ob�fd Ԟ2��,& X�OCA1E!��$OP����V�t ����P��Pd��`RŃ�aOUx��3e��R�5Ie h|�1��e$PWRL�3IM;e�BR_�S�40��� �3H1UD���t�QBte7�$HSu�!�`ADDR2�HB}!G�2�a�a�ac��R��x�f H!�S ���u��u
�u��SEv��"�HySH�:g $����P_D�H Y�RrP�RM_����HT�TP_i�Hx�h (*�OBJ���b��[$2�LE�3�s>�i � #�"��AB_
�Tp#�rS��Px���KRL{iH_ITCOUw�B6�L`�rQ��U�`̹�`SS��JQ�UERY_FLADQ1�pWR�N1x�jp�gP��PU����O ���q�!t��/t��~� �IOLNw��k(�� CJq$�SLL$INP7UT_Y$;`���P,��̀SLA.� l׀�(�`$��C���B��IOgp�F_AShm}��$L��w��8AِU � 4@_1��݃��情@�HY1ǧ�����[�U;OPen `l�ő�2��������[`P �c;`�	������2}Ja�o � K�CNEaG4�v7F�Da�֏2J7VpOQR$+J8q�7�I_1z�>��7_LAB�1�Px|���p�APHI���Q{���D�J7�J�-��_KEY�� �K��L�MONx�p�$�XR_���)�WAT�CH_��C��D�E�LD��y�P��eq� @Р1V�@&�U�C�TR�3U�i����L}G��r� !#�LG�Z�RࢵcX��c���FD��I�� ��\!����� ����e� Dqf�ce�c�e�ΰe�@� e���@0J_�� �1j��qʦ�F�Ax�ȒĞ�Cd(��SB����c��c���ΰ��I�����ƍ ��枰RS��0  M(w�LNe�<sѐ���)��6Ѽ��UosD��PLM�C�DAUi�EAwp���T��u�GH�R�ao�B�OOw�t� C���`IT\���� ������SCR���㇑�DI��Sw0HRG X ���z�d(��o���w�W�o�X�z��JGM^�MNCHLl�n�FN�a�K��7PRG��UF��B�n��FWD��HL��STP��V�� ��,�Г�RS�HzP��w�CdD��1Rz�: :�^�Unq��9���H�k�����Gw�@( w���0����s�}�OC/ ��EXv�TUI��I��7�C�O�`����<@���	$���<@��NOANA8o�A2� VAI���t�CLUDCS_CHI$�!s�O�L
�SI��S��IGN���ɳ��rh�Tc�DEV<�cLL�Aʀo�BUI ��uP�j@T��$��EMr���]�.+!	1vP�j@ހ���~p����1�2�3����� 
0w ��C��x�Q@5������IDXa$9 [����֥1V�STƐR��Y}��<@   v$E.&C.+�pmp=&P&�!��	1x L����`���4@r�`Na�eEN�wp�d/�@���_ y ap7�}p	b����#�MC7�z{ �C�CLDPƐ>UTRQLI��T8T�94FLG)"0��Q53�DD�57t�LqD55455ORGT� 8�H2_ȲF�8!s�D/r� �#�S{ � �	59�455S�PTD0��0y0�4�6RCLMCD�?�?Iƀ�1�PM�p^����|�$DEBUyGGugQDATAY�r�T �UFE���T)!�0I6p�T} Yd@��RQ��0ODSTB�`� V��D��HAXR��G>�LEXCES$R�aR�BMZ`��~��B�4�2�ASq�����F_z@�H�S[�O�H���MJPTH��� &Pv�m��QMI>R� � � [w]R�RCT��UN}��VO�ZA�ZL�RC�PC��Q�`�D��O�^�CU_RPX_THqG�P�`R`|1��)`/d55�R^`�`S�P �B_�FR@^�a\fZ_���^ddpG��* �w�MKH�� \���r�Fv$MBu�LI��q�cREQUIR-EG�MO�lO�kfB�Kq�ML� MG�� ap���`|��cB]i MNDU�Sz!�>�5�Z�9sD��Q��IN�p��Q�RSMPf�Sx� �Q�!E]�q��&rPST� o� 4�LO�Pf�RI ��EX�v�ANG��A2�1�A5QG���@$�QG��MFh������"���%&�2ТfSUP��%�!F `RIGG>�� � ��0�#�1��Ӫ#Q��$$���% #n�א~�א��rP��8wAZw@ETI9���12�M\p9� tV�pMD�I��)��� �DA�H�pu���DIA���ANSAW,��w���D���)�AO7��0�Љ �QU��VB�70�vr�_V@�ъ �C�0��sX@�b|ٰ���P���v���P��KqES�!���-$B����� ND2FB���2_TX�$XTR�A�1����`LOāЪЋ$RG��B�F�8Ҍ|�g�_��RR�R2�E�0 #�W�e�A�1 d$OCALI�@2�G�:��2�RIN����w<$R��SW0"D�ᣫABC�xD_�J��a����_J3:�
�1SPs�rp��P�-�3,���?�
��\�J�l��2�1�O8IM� �2CS�KP":��~�YÛ�J���2Q��̵��̵·��p_AZ�2h���E�Lg�FAOCMP0�s�1!I�RT�A)��Y�1�i�G��1��K�> Y�ZW�SMG��܀�4JG� SCyLP�uSPH_� ��0���������R�TERࠧ���[IN��ACz�|�`�� ��r��} _N���������1i ��?R�� �DI��0�pD�HP3��ё�$aV��Rs��>$v� �p�1������E��H �$BE�L�?w��_ACCEL��ث���PS_Rـ0�QT!Z�*aEX2L6b ��3���׀c��.a��h���36cRO
Q_�m�J�P��2�p`��_MG�$D�Dm�����$FW��0݀�Ӊ�Ӥ�~�D}E��PPABN��RO��EE`���0±�YAOP��6`Ra_��YPaPC��YY����1 �!YN�@A��7����7�aM�A��ig�OL�de�INCa��q�����B�����AENCS���Á�B�Ѥ��D+`I�N"I6b��ހ��N�TVEk���23�_U�����LOWL�#F�0��DF�D�`��� ��`R9C����MOS� wT�PP�2��3PERC�H  8OO`��  z�q�!�4!$ǐ�!�)b��A6b�L �tW����F�
�4TRK��!AY [�(cOQI6bXM�pp/�SQ�� MOMc���BOR�0���D�㣧0d��⍠DU��7b�S_BCKLSH_C6b��@YO`?�������*N�ĵCLALM���1�?P6%�CHK0� �GLRTY������Ѕ|1r܁_�N_UMzC��&CzC{���#��LMT)�_L�0ú$+��'E�-� �+� �Հ�%��>��C�!4�P	C��HI��`q�%�C@8�{��CN_b��N"C�6��SF���	V!�p!����U16b��5Y8CAT�.SH �����?a���X�07aX�L�n�PA�$��_P�%s_����P n ��`rDc%JAaP�fC	 OGs7�TORQU�A�Li��`�bd����B_W� IU�n��D_��Ee��EUI�KI[Ie�F�P`�As�JX��w�VC��0�jS1q^o��_��wVJRKq\�R�V�DB��M��M�Pp_DL_��GR�V�D�T_��Te��QH�_^��S�#jCOS0k1�0hLN�PSktU Zd_�Uiv�Ui'Q�jl�EQ�UZN`d�QMY�\a�h<b��Dk�iTH�ET0$NK23�e�rY�]`CBvC5BY�C��ASrqDr`'TRq_�RqvSB_Ӝpr*uGTSֱ��C�0��qO�;C_Ǧz�c$DU` ��r����xR�v���Q��53�NE��7�I^`q#;��$=�qAu;�D�8"e-h-aLPH0e����StU��e���e@��f�����f=�V]�QVR�O�u�V��V��UV��V��V��VɋV׉H]���|�t��1T����H��H��H��UHɋH׉ON�O]��O�s�O��O��O���O��O��OɋO�fF�?q��e��P��SPBALANC�Ec�=1LE�pH_uSP��pf�f�>�fPFULC�������e��1�+�U�TO_[ �ET1T2_���2NB!���� ����� ��p�ҚӞ�T
O����@IN�SEG��=REV8��= ��DIF3ٳ1��1�1�&O!B�&!�S�2�@���M!�TLCHWAR���&�ABBA�$MECHHq�`V�\�q&AXVP4u�4�@�T�� 
v��Ab�n��ROBn CRyB���j2 �MS�K_֠�ԓ P j�_�R���2����51�2���������$��>�INű�MTCOM_C\P>�Д  h��~��$NORE���Q��.�@�� 4�@GR�Ba�FLA�ű$XYZ_D�AQ����DEBUb�� f�.�mЖ ��$/�COD! ��҇b��$BUFINDX��w���MOR��� H�����E&���~�^�$޲��1o1�� TA������аG�Ҙ � $SIMULp@�С��\��OBJ�E��\�ADJUS<z�m�AY_I�A�D��OUT�@�Ԡn_�_FIb�=��T�@��������q���������D,�F�RI��T�RO�@��E�A�OPsWO�P���,�ПSYSBU+���$�SOPT���;!_�U<^��PRUN0҅�PA��D��`�Y� a_��2z��AB���
0��IMAG!4���PϱIM����IN�P����RGO�VRD�v�e��P0����� ��L_R�zA�(�"�0RB� � >1MC_ED��b� 
0N+�MW	1��MY191  ��SL����� �ޡ�OVSL��SDI5�DEX�3��3$
�V�@�N��A���� ���n�Cb�0T����{�_SET�@��� a@�@!��RI^���7_Lq@YL� 	���x�0 ����Ta��@AT�US�$TRCp���ҔBTM��I��l41sU .��� D��E���4�E���� & �EXE�r!L�� "�)�0���U�P��!IS��X�NN��1ldQ���PG>՟L�$SUB��V�Z�JMPWAI�0P��%LO� ��̰[��$RCVFAIGL_C�i�!R�� i�r�e1�0�4���%�`�R_PLZDBTqB�A�2i�BWD�&fY�UM�@�$IG��8�����0TNL�0�$@2R'�T�~@�@��P�PEED5 �3HA�DOW�@c�Y�f�E��4�p!DEFS}P�� � L���|��0_�0���3UN!I����0C!R �L�`̰P�5�P1�����Ю@^Ѻ�� ���N�KET�B�@��AP42���� h �pSIZAEy@������`ASx��ORZFORMATK�*4CO~ \Aǲ�EMn�|D�3UX8C����PLI%2���� $I�OMP_�SWI/��E��W4i�Js��AX
0%0?AL_ ��@�0�"�gPBJDpC�D��$E!�J�3D�H� TV@P�DCKC m�CO_J3r�RQRĢ�l	_] ��@C_/1�A  � �h�PcAY�qҧT_1�Z2�S�@J3�p�[�Ux�V�S6�TIA4�Yu5�Y6�MOM�@c$cc$cc;�B� �ADcHfcHfcPUSpNR)duecue�bx�B�ħ` I$PI��U���U *s�Uus�Ujs�UUt�f �kit�t��v��v_!���m���:v3HIG�Cv3�%�4iv�4�% � ��iv�sxx�!�y�!�%SAM����tiw��s�%MOV��$� '�
�ް)p%��� #� �0�P2��P%�0�5�`�!��@��H��#�IN j��@�sq���h��"s�𳈊���ӋGAMM�Ǧ���$GETH���Є�D�T/�
z�OLIBR9!W2I��$HI8 _��%�H�E"�U�AO�r�c�LWJ�����r���c��Rn�M0�AC50� �a ?^I_ �p2�/��B�X�AY���$c/�Hf��C {�$,X 1���IXRk�D�>�A!�$@�LE ���`����Xq��Z0MSWFuL�$M�@SCRI(A7���)q�T"��C�����P��UR��$�v�KS_SA�VE_D-B�;#NO�PC`<"�TB�&� �_�a�YW��i�Y�`��@��pkR#uܸ�SD�� �p#�s0�@�,�$�cx Y�sv�x@�<�����<!BL���ĩ � "�YL�c��Y��S��6�0�� 0 ����J��������	�t�Wq����`��d1�t�M����CL�Ȑ�Q��o �1T"�@M�3�*� � $��G$WRГ� ���QR�oTP�vTP�}T P�T0���+��C;J�@X�0O~S�AZ�ո�@��Uԫ �ՑOMK��V��������̿`CON�� �A�PL�Q_v"� | =Q�B�$i��c��c B��Z���j�A ��@(�P~����@�P���P_A�PM� QU��p � 8@Q�COUM�i�QTH�/0HO��G�HYSf�@ES�F�UE2�t8�@O�D�  �@1P0�@�`UN�����t�Vr�а P�����%$��W2RO�GRA���2�O�����IT����t�IwNFOXѱ �Ah������OI�� ((�SLEQ@Zv/Nu/ ��+S���s$� 4@EN�AB~�� PTIO�NZ�4(r��4cG+CFl�0J� �AV���,�R��|�BOS_ED� N�е �N��K�j:G�E��NU�AUT^�CO�PY�8 7�1j�M�N�NAE�PRU�Tf� HN� OU��BN�RGADJ�XѶTBX_t��2�$�0��мW�P�����v3��#EX�� YC~���RG�NSh���ޠLG�O��PNYQ_FREQ�bW��MvM!�D��LA��D!�c��@CRE3�R����IF�a��NA�q�%�$_G}4TATxB0�$>�MAIL�r 2��!��B��1�!1�$�ELEMl� �|s0vFEASIy @��L���2@K�66�V�2�I��0�D"Eq0J��k2AB�AP�E��vpV�!�6BA!S&R�52��aU�p���W�$�1�7RMS_TRe3�A���3 �ӓp�r�!�4�B!"������	B2 2� ���ԇ�(F�2 'G�2/�_����2SG�gN��DOU��N��!"PRe�m �6G�RID��b�BAR�SZwTYz�U�O\?`Xѻ ��_�$�!��B�DO��i�� � ����PO�R���C�f�BSRV�� )TVDI`�T��P0QCT� MWCpMW4�KY5KY6KY7KY8�/QM�F�l��$VALU�35�(4�2��Qi��C uY����C�!�2�� AN4��R�!R�R!2�TOTALX�s�a2cPW:#I�A>HdREGENFj[b��X�8��R%��V-�cTR�3�rFa_S8��g[`�V���b��2E�#�@L�1�-ncV_H�@DA-��`pS_Yf���^&�S�AR-�2� }�IG_SEC�ȴ`R�%_���dC_�F�Q�E�q�OG6�kNjxSLGEpl�� �>�_%��/�0`9`S,���$DE.QU>���̧�pTE���P�G� !�a��aJ�v<^�3IL_Mm$;����`��TQ-�6���0Ƨ��Vh�Cv�Ph�#1��M��V1���V1��2��2��3*��3��4��4��$���`ӓ%�� 0����INA�VIB=�p�]�T�d�2`�2l�3`�3l�4`�4l�X�WB���SB����D ?$MC_FP���%�LC�B�f#c�Mo�I��oC ��6��qL�KEEP_HNADDᑑ!#��0-�C�ѫ  C��A⒤�D�O&�"��{��3�D��!a#D�REM[�C�8a�B��ԗ���U�$eC�HP�WD  #�S�BMSK�BCOLLAB/��P@�$a�" IT$ ��fȕn��� ,(�FL{�LW�M�YNڐ1�M���C`r�G`UP_D�LYX���DEL�Ac�9a�"Y�AD�-�q�QSKIPNw�� �P��O��cNT9�����P_�� ����ҏ�÷�aѹ �ѹdPкqPк~Pк@�Pк�Pк�Pк9�O�J2R ���qX�0TG#r���qr��� �r����* RD]CS�� �_�R�R1�o�I�R�!��J���*DRGE� T3���BFLG'����*D�SPC��!UM_|r�!�2TH2NrA�<�e� 1� g��@� 11��� l����O�v�ATy��.��Q&�� W ���� *D�Ҙ�I��H��ҥV�2]���c�u߇ߙ߽߫� U�3]�������X�(�:� T�4]��]�o�������5]���������"�4���6]��W�i�{�������� U�7]��������
.W 	U�8]��Q�cu��� U�S|�L�  �1�V�p`�W���E%$�рp�e)fcI�O��Ip��R���WEC�� �M0���!i�$c y�+��$DSB] �� �""c^�CB�p�� <M
E�+��	D���0E�"��MDt"'��M�E� D�p^�'DBG_~@PD��3%!eaPG
A@�x��R�S232i'� ����P��pICEU�2!`k$�p�ARITq!aOPyB�rFLOW>p�TR(.b��@qC�U� M%3UXTA��qINTERF�AC�$��U`���� CHA׃ t�ݐ"!hp��$�`�`OM'p�sAD���0Iᓴ0Q@A+��TDSv`���8c3�EFA����r�S� k��`8b� q��R H��6A �ٶ�q  2�� �S��M �	O� �$)�s�0��
eC2`_%pFDSP)FJOG�`�#�p3_P���"ONg�u���'�	6Ky0_MI1REAb$wpMTY��CAPK�wp4Ц@�4"A�Sp}@r"At �EBRKH<16=��R��! �B�s�BBPo0�b< C@BSOCF��uNUD1pY16���$SVi�DE_�OPGtFSPD_�OVR�k��DLTRWCORbW� N�PbcVF�@�WB@OVEECSF�Z^p�S,rF�V� t'�UFRA�ZTO�$LCHa�u�2�#OVST��B@WQ����BCZ� r&PQ@]s ; @�TIN�``!_$OFSC`C�0@�WD|QdxQ%Q�,�E?PTR�!e"�A�FD���AMB_C��bB5@B<��!q�b�a�cSV��L�k0ȉ�s��RG�g�HAM�tB_=0�e-b_�M�`2�:`T$SCA8@�D�B?p�HBKo1~6TqIO��cu�pqPPA Wz�qhy�t{uu�:bDVC_W R#�p1 ��p���Q�u���x-s�u3�v3`��{�0p@�SQUR#7@~CAB ���,Ӟ`���`�h9��O�`UX~6SUB'CPU�O@S��� ���dp0ݱ���c�d�~��$HW_C]� �0ݱrpʆ�� �NÐ�$U��D��>�ATTRI�0���O@CYCLw�NE�CA)��CFLTR_2_FI�/����LP[KCHK�ՠ_SCT�CF_��F_�|��FS8��b�CHA��d�p���b�"��RSDU�`�Q�3��_T�h0Y���c� EM"��EM�CT��ݰĀ�����2�DIAG5R�AILAC�sx�M���LO	P7�/V����3� H�3��sPR��pS+� 90��C��q&0	,cFUNC:��1RIN���a$D����!ʰS_"@*?p䣸�Mt����MtCBLȰ���A0�
��
�DA�@�O���LD`0GPpq�w�*A�|�w�TI�����AĀ$CE�_RIA��AF�Pn#ò%`ȵT2bd�C}3�r�aOI��fDF_LY�Rl1��0LM`#FA  H�RDYO�AM`RG�|�Hސ�Q� W��MULSE��3��8P.�$J_ZJzR�W��[FAN_ALMsLV�#��WRN��HARD�@o6���2$SHADOW  `������V���!�Q��E_`s�AU��R���2TO_SBR ��6@(�逺sá@�_MPINF8`��8S�m�^�REG���DGy�K�Vm0��F�DAL_N�dFLۅ9�$Mm�l��hg O`L�K$g$Y("V1��2~#�� ��CCEG[ CGP
�A �~/U28S�;��EA�XE,GROB)JR�ED)FWR  �A_i�SSY�@D��@��S��WRI  �ɀ�ST�*C0�@nPE��&�w� �"@B���9a��5k�pOT�On�%`ARY�)C�e����[@FI��@pC$LINK��GTH2��0T)_��9a%�69R[�XYZo2e�7s�OFFA`2� \�N�uOB'@����a� h0��FI���0�4?T��AD_J�!�2@lR?�pq������89R � ��	T�AC��F�DUWb$�9x�TU�R��X��z!�N�X��� )FL[��PH�0�� |���309ROa� 1�KN@Ms�/U3��{�������W3ORQ�6A��(��{��@O��N��Hp�34A��]OVEd("M00J��~��~ ��}F1|J�|�{AN��5�~ȱ)!e }@���ve�%0��%�6AERSA	|�E �`��E$A�Ā��ܥ��V�S�V�AXc�2V�� ҁ4�%8��)b��)w� �*�*r�*��*: �*q �*1� �&��) ��)��)��)��) ��)�9�9�'9�D189DEBU���$����<��1VbV�A!BV�Tq|Q^VIp�� 
B�s��+E�� 7G8Q7Gw�7G�7Gr� 7G��7G:7GqδF �Ȳ4��LAB��8)���sGROB�)��2pB_�,&�� uS��%��FQ*U�VAND� |�:$3�_�=!�YW 2qZ�^�`mX�|X5�^�NT��
c�PVEL���Q�T��V�SERVE��P��� $���A6�Q!�PPOHb����`��Q�R�����  $bT�RQK�
 ct�
`ߌgȲ2�e��Q�_ � l���a��'ERR��m"I� �P��raTOQ��L�H�$��f�G�U%�H�f�   c��	a� ,�Q#e=`��R�A�a 2� d��b{s�Ta ���$r����"� cOCG�p� � dkCOUN�T�� �SFZN_CFG	aG� 4ƀ��;�T�� ����3����m!�pRs^��� �(@M���o���#������uF!A���ö�sXd��{ �y�a��S��TO�d�9PJ���HEL��Yr�� 5k�B�_BASf�RSR�֤�^�S끐�M��1�gM�2p�3p�4�p�5p�6p�7p�8�g@�ROO��`9�f]�NL��LAB�S�N�N�ACKFIN2pTo���$U��M��� �_PUV���b�OU�P̠��-��f������&TPFWD�_KARwa��f`R�E�T,�P/�]��QUE���eU �����I��C-�[�[��Py�[�SEM3A�AA�H�A�qSTY�SOސ	�DI�ɠ}s����'��_TM��M�ANRQL�[�EN�DZ$KEYSWITCH^�s�.��ĔHEU BEATmM��PE�LEvb(��@��Ur�F�s��S3�DO_HOM�ưO���EFA PAR��rv����C���O8�c`�aOV_Mx����IOCMGd˗?��.�HK��G� DX�׍pU��¹�M����HFO;RC��WAR(�	��,�OM� � Q@�4���U��P3�U1��2��3��4=�V�@�SpO��L��y��b��UNLO9�����ED��  ~�PNPX_ASZr�� 0�ЄЍp���$SIZ��$V�AP�eMULTI�P��.�ŰA��?� � $H�/�H���B�S}s�Cr`���FRIFm"pS���������NFO�ODBU��~P������>�UD_Y�SN��з� xU`SI�bTqE�8��SGL*�	TA� &opC��C���+�STMT�\�P���BWe,�SHsOWd�n �SV7 �_G�r� : $PaC�@p7#�!FB��-P��SPːA����"pVD�Оr�w� �WaA00^T ��ɰ��Ӱ��ݰ��簪��5��6��7��8*��9��A��B�ٴ� �׳A��y���F��70T���1�1"�1/�U1<�1I�1V�1c�U1p�1}�1��1��U1��1��1��2��U2�2�2"�2/�2<�2I�2V�9 ���p�2}�2��2��2
��2��2��� `�>`"�3/�3<�3�I�3V�3c�3p�3�}�3��3��3��3���3��4k	4�4��4"�4/�4<�4�I�4V�4c�4p�4�}�4��4��4��4���4��5k	5�5��5"�5/�5<�5�I�5V�5c�5p�5�}�5��5��5��5���5��6k	6�6��6"�6/�6<�6�I�6V�6c�6p�6�}�6��6��6��6���6��7k	7�7��7"�7/�7<�7�I�7V�7c�7p�7�}�7��7��7��7���7��)�VP��Ub� `{@e�Q
�����Q�U�PMR��CM�p�bM�P�R9` ��TQ_+pR��P�e(a~��Sn�YS�L�`�P� �  L��jw��A�ؠ; Ѡ<�D��VALUju%��x��A6XF�AID_YL��^UHIYZI��?$FILE_L��T�i�$��P�CSA~q� h �pVE_BLCK����RE��XD_CPU �YM��YA�us�_�TB`�Y*�F�R � � PW-p��6<aLAj�SqAc�RaKdRUN_FLGde@dhaKdv�ke�a@d�aKeHF�Wd�`Kd�� 
�TBC2��u� � �B k`(���pĠ���d	�'TDCk`|r�b�p��
u�gTH	�%s�D�1vR��ESERCVE��Rt	�Rt3����`�'p �Xw -$}qLEN��0�t	�}p)�RA���sOLOW_�Ac1}q�vT2�wMO�Q�S���I.��B�Q�y�D�}p�DE���LA3CE,��CCC��B��_MA2��J� ��J�TCVQ�r� �T X�s���������Ѷ�$ ���J+���Mۄ~��Jw������ ��q2��������JK(�VK��:�>��:�sq/�J0O�>�J�JF�JJN�AAL�>�t�F�t�n�4o�5/sX�N1����d�N�
�DL�p_Xќ�uA�`�CF6�� `�PG�ROUDPF�Q���N��`C�� �REQUsIR=rؠEBU���yq܆$T�2��6�zp ��$$CL�AF� ���4Z�*�*� O����X�e���~k�IRTUALW��i�AAVM_WR�K 2 ��� 0  G�5a�ͯ٨ʯ.�� ��	s@�3�*����!�^�E�c���������ɿۿ�㴧�BS�@�� 1�x�� <��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<�~pN�gLMTu�?��7  dQINZl�PPRE_EXEb}� �~AAT��ʖ���IOCNV�Ւ~ �hP�UqS���IO_� w 1��P $����I�4��1��?� ?_ Tfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο�����(�:�Q L�ARMRECOV� �c�L�MDG �(BLM_IF m?����� �+���N�`�r߄ߕ�?, 
 �߾߀9�E�������A�NGTOL  ��
 	 A  � Y�k�Q PPLI�CATION ?��� ����ArcTool� �� 
V9.?00P/03j�+�
88340�����F0����161�2�������7D�C3��+��Non}e+�FRA+�� 6�LP_�ACTIV�	�j��UTOMO�D� �Ո	P_CHGAPONL��� ��OUPLE�D 1� � !3��CUR�EQ 1  UT=	==	�������=_�ARC We=l=�AW�ՕAWTOPK�HKY�Dy�9 'EK]o� �����5/�/ #/A/G/Y/k/}/�/�/ �/�/�/1?�/??=? C?U?g?y?�?�?�?�? �?-O�?	OO9O?OQO cOuO�O�O�O�O�O)_ �O__5_;_M___q_ �_�_�_�_�_%o�_o o1o7oIo[omoo�o �o�o�o!�o�o- 3EWi{��� �����)�/�A� S�e�w���������� ����%�+�=�O�a� s����������ߟ� �!�'�9�K�]�o�����OTOC�����DO_CLEAN��|���NM  H���^�p�������A�_DSPDRYRL���HI��<�@M� �&�8�J�\�nπϒ���϶������ψ�MA�X��������
�X��������PLU�GG����
�PRUC˰B:�H�����d�Oi�Կ��SEGF��� ������:� L��&�8�J�\����LAP������ ���������"�4�F��X�j�|�q�TOTA�L,�U�USENU
���� ߨ���O �RGDISPMM�C� ��C���@@M��O���߹RG_STRI�NG 1��
��M��S���
__ITEM1i  n����� ����'9 K]o�������I/O S�IGNALc�Tryout m�odejInp� Simulat{ednOut-,OVERR = 100mIn cycl!%�nProg A�bor7#n$s�tatus�${ c�ess Faul�t�,Aler�$	�Heartbea��#�Hand Broke���/?�?%?7?I?[?m??��e��w�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O__�?WOR��eKQ �?%_s_�_�_�_�_�_ �_�_oo'o9oKo]o�oo�o�o�o�o�nPOc�!�`c[�o$ 6HZl~��� ����� �2�D�8V�h��bDEV�n�� ����̏ޏ���� &�8�J�\�n����������ȟڟ����PALT�=7�c_�_� q���������˯ݯ� ��%�7�I�[�m��8����%�GRI�e ۱O�����'�9�K� ]�oρϓϥϷ����� �����#�5�G�ɿ��R�=��Yߧ߹��� ������%�7�I�[� m�����������m�PREG;�$�� ��K�]�o��������� ��������#5G�Yk}���$A�RG_KPD ?	�������  	]$�	[�]����� SBN_?CONFIG� ��%!$"CII�_SAVE  ��D;� TCE�LLSETUP �
�
%  OM�E_IO��%MOV_H����REP����UT_OBACKs�	�AFRA:\�� ��^'�`� �<(� �M+@ 2�3/04/01 �14:33:48���/�/�/�/-,��?/?A?S?e?w?�?��?�?�?�? �?�?O�?5OGOYOkO }O�O�O,O�O�O�O�O __�OC_U_g_y_�_�_�_�Ё�_�_�_�_�oo1o�OINI�:�o%7#MESSAGS]a^� >hkODE_D�V�7G�eO���o#P�AUS�a!��� ,,		�� ��ow�o- 9;M�q���������;�����d�`TSK  ��m</Bo UPDT̖`[gd���fXW?ZD_ENB[d3��STAZe�����WEPLSCH �R+   b��.�@�R�d�v� ��������П���� �*�<�N�`�r����������̯ޯ����R�ODނ2��4���/��>� % V�{�������ÿտ翀����/�A�SϾWEROBGRP`���r�GWEWEL �2�D���h��� ��'�9�K�]�o߁���ߥ߷��߼	XIS%UN���D��� 	r����@� +�d�O��s���������METER 92b�_ P��&����J���SCRDC�FG 1�N! �[[?� ������������5/�
QW��M_q�� ��2�%�7I���!GR��Р��o�UP_N�AME 	��	�$�_EDY`1�s�� 
 �%�-BCKEDTA-v��/*/j��  �����.��µϰ����/:����%2 �/���/a/��G(�//? v/�/?�/�#3g?�/ �?�/>�?�?B?T?�?x?�#43O�?�O�?>�\O�OO O�ODO�#5 �OoOL_�O>(_�_�O�O�__�#6�_;_o __>�__o�_�_No�_�#7�oo�o+o>�o@+ro�o�o�#8c/�//�=��>P�t�#9/��|���=X�Ï
����@��!CR�/�oG�Y� }"���ԏ�|�
��~�NO_DEL���GE_UNUS�E��IGALL�OW 1�� �  (*SY�STEM*��	$SERV_u�.�G��POSREGP�q$r�.�G�NUMu�<����PMU����LAY��.�PMPALTǧ�CYC10Ԟ�xѠծ�ULSUǯ0���r���L#�\��BOXORIy�C�UR_I���PM�CNVæI�1�0����T4DLI�B@�b�	*PRO�GRAO�PG�_MIծ���AL(ߵ���B<�G��$FLUI_R�ESU�u��j�������������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r�������������e��LA�L_OUT �6�q#�WD_AB�OR��i�ITR_RTN  �����l�NONST�O��� ��CC�G_CONFIG �7�7���8������E_RIA3_I���, ����FCFG �����5_L�IM^�2� �� 	n���Q<j�ߥ蜀�d�PAV�GP 1.?���-?�C�� C_�  C�b�fU�b�f�f�b��f0�D`�DDU��
��i���Dv�DZ�l~�����x�D/�9�C��M�W�a��?���HE��u�"�G_P��1� ��d/v/�/�/�/�/�/HKPA�USf�16�, ���/ ?6�?L?2? \?�?h?�?�?�?�?�? �?O�?6OHO.OlO
�O9?��h�COLLECT_9as	`�N�GEN߰p��~��B�ANDE�C�s���1�234567890!W��a�O_1V��'
 H+���)l_�_ a�k_}_�_b��_�_o �_�_	obo-o?oQo�o uo�o�o�o�o�o�o: )�M_q��������Fm��K �N�FIO !
Y�A�����������ʏb�TR� 2%"F�(��}�
�؎���#q�� %[�_�MORm$� � )���������ǟ����ٛd��n%r�,� %?	!	!�>���KTH���$R9&�O�w�v�v�C4  A���
� x��A>A�Cz  B�fP�B���C  @֘������:d��
\�IS'f��\�T_DEF*� ��%�+�����I�NUS�&,@�K�EY_TBL  ��,v� �	
��� !"�#$%&'()*�+,-./*W:;�<=>?@ABC��GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾��������͓��������������������������������������������������?������6�d��LCKI���d�I�S�TAs�>�_AUT/O_DO��m����IND�D�δAR_3T1�Ͽ�T2���ز���A�XC� 2�(q�cP8
SO�NY XC-56�{�u��U��@����� ��А;~�HR5XY ���߭�R57����A�ff���6�H�  $�m��Z������ �����!���E�W�2��{����TRL�L�ETE!��T_�SCREEN ��
kcsc�"UD�MMENU� 1)�	  <u��1�: o`CLr���� ��� &_6 H�l~���� /��I/ /2//V/ h/�/�/�/�/�/�/�/ 3?
??B?{?R?d?�? �?�?�?�?�?�?/OO OeO<ONO�OrO�O�O �O�O�O_�O_O_&_ 8_^_�_n_�_�_�_�_ o�_�_oKo"o4o�o Xojo�o�o�o�o�o�o��o5+���_MANgUALH��DB9��0�����DBG_E7RRL�*����� >���~~uqNUMLIM�����dn�ޠDBP�XWORK 1+���L�^�p�������DBTB_�� �,�}����u��RqDB_AWAYz}s͡GCP n��=����_AL
����yrYGл�n��nx_�p 1-q�́.�
;�y�z��g�����_M��IS����@A���ONT�IM���n���ޖ4�
X�I�MOT�NENDM�H�RECORD 13��� �����G�O�t�b���������į ֯m�ޯ�t�)���M� _�q������˿:� ���%���Iϸ�m� ܿ�ϣϵ���6���Z� �~�3�E�W�i��ύ� �ϱ� ��������z� /��:���w���� ���@���d��+�=��O���s�^�l�����Oi������b�8M��sN��������[���);�_J8X���W�����N/��9/�k�0.:/q/�/���TOLERENC��sB�>��L��up�CSS_CNST_CY 24,���p	�/<���/??(? >?L?^?p?�?�?�?�? �?�?�? OO$O6OHO��$DEVICE ;25�+ І�O �O�O�O�O�O__+_�=_O_���#HNDG�D 6�+ՀCz�i^LS 27�M a_�_�_�_oo'o9o�c_�"PARAM C8U�%�duKd�$�SLAVE 9��]nW_CFG �:koKcdMC�:\� L%04dO.CSVJo<�c�olfr+"A sCHp��Q��Kn*_}g�KfOr|q�zyyq�`JPѬsk~<�ρ��lRC_OUT� ;�MρOo_SGN <K�4��a�01-APR�-23 14:3�5p+�=��F V�t�g�c�Knd����mE@�S�Þ�j�x��z��cVERSIO�N �V�4.0.1��EF�LOGIC 1=^�+ 	�x�`���q��PROG�_ENB)��V2�U�LS� �V�_�ACCLIM����c�q�WRSTJNɐ�3��a��MO;�uq�b��I?NIT >�*K�v�a ��OPT�`� ?	�Ȓ
 ?	R575Kc��74!�6"�7"�50F�ׄL�2"��xp�|އ��TO  ��z�ů߆V֐DEXҞ�d���pݣPA�TH A�A�\˯*�<��+HCP�_CLNTID y?�c �{�G#|��!IAG_G�RP 2C�i Q�	��ؿÿ���� ��Dϒ�m�p1m10 89�012345678n���=�� ?Ϝ� �ω������r��� ���!�3���\�n����q�Gߩ߻ߙ��� ��{����9�K�)�o� ���U�g�������� �����3�Y�7�i��� �+�u������� ��/gyW�� 9���	�-? �>χ:ϫ�� ��|���;/&/_/�˰_O 4Q/�/A/ #�/g�/?!?혒$ -?W?�/g?�?o?�?�? m�?E/O�?ODO/O hOSO�OwO�O�O�O�O��O
_�O.__R_��<�p c_�_�_ C_�_�_�_�_�_o0o �_@ofoQo�ouo�o�o��o��CT_CON�FIG D��|ʓ]�eg�u���STBF_TTS��
J�)s��}�xq:<v�pMAU��?�~Q�MSW_CF�`�E��  ��OCoVIEWPpF�}�a�������� *�<����e�w����� ����N������+� =�̏a�s��������� ͟\����'�9�K� ڟo���������ɯX� ����#�5�G�Y�� }�������ſ׿f������1�C�Uϡ|RC�sG]r!�c΍� �ϱ�����
���.�t�SBL_FAUL�T H�ʥxH�G�PMSK2w[��`TDIAG Iy�qUt��UD�1: 6789012345��x��c�P�o����*�<� N�`�r�������@������;�Vp����@8r��\��fTRECP�ߣ�
�ԣ��� ��������1C Ugy��������	0�B�?f�U�MP_OPTIO1N2pT�aTR�r3s:X��PME1uu�Y_TEMP  È�3B�Vp���A��UNI�np4u���YN_B�RK J��bE�DIT_y�ENT� 1K��  ,&�R/P@/}/P�l/�/�/�/�/�/ ?�/'??K?]?D?�? h?�?�?�?�?�?�?�? �?5OOYO@OhO�OvO �O�O�O�O�O_�O1_�C_*_g_N_�_r_ MGDI_STA�ؔq�%NC�S1L�{ ��_�_P
Pd7Yoko}o�o �o�o�o�o�o�o 1CUgy��� ������ �.� Fa.�T�f�x������� ��ҏ�����,�>� P�b�t���������6� �����#�=�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������۟���	� �5�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ӿ������-�#�I� [�m��������� �����!�3�E�W�i� {��������������� ��7�ASew� ������ +=Oas��� ������///9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?��?�? �?O'/1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�?�_�_�_oOo ;oMo_oqo�o�o�o�o �o�o�o%7I [m���_�� ��o)o3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ����џ����!� +�=�O�a�s������� ��ͯ߯���'�9� K�]�o��������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߷���������� �-�?�Q�c�u��� �����������)� ;�M�_�q������ߝ� ������	���%7I [m����� ��!3EWi {��������� ///A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�� �?�?�?�?/O'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�?�_�_�_�_ Ooo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu��_ �����_��)� ;�M�_�q��������� ˏݏ���%�7�I� [�m�������ǟٟ ���!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ� ����������'�9� K�]�o�鿛��߷��� �������#�5�G�Y� k�}���������� ����1�C�U�g�y� �ߝ�����������	 -?Qcu�� �����) ;M_q��y�� ����//%/7/I/ [/m//�/�/�/�/�/ �/�/?!?3?E?W?i? ���?�?�?y?��? OO/OAOSOeOwO�O �O�O�O�O�O�O__ +_=_O_a_{?�?�_�_ �_�_�?�_oo'o9o Ko]ooo�o�o�o�o�o �o�o�o#5GY k�_�����_� ���1�C�U�g�y� ��������ӏ���	� �-�?�Q�c�}���� �����ɟ���)� ;�M�_�q��������� ˯ݯ���%�7�I� [�u�g�������ϟ� ����!�3�E�W�i� {ύϟϱ��������� ��/�A�S�m���� �߭߿�ٿ������ +�=�O�a�s���� ����������'�9� K���w߁��������� ������#5GY k}������ �1CUo�y ��������	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?gU?�?�?�?� �?�?�?OO%O7OIO [OmOO�O�O�O�O�O��O�O_!_3_E__? ��$ENETMO�DE 1M�5�  o0�o0j5�_�[nPR�ROR_PROG %{Z%i6�_�Y��UTABLE  {[�?-o?oQo_g��RSEV_NUM� �R  ���Q�`�Q_AUT�O_ENB  ��U�S�T_NO�a �N{[�Q�b W *��`��`��`	��`�`+�`�o�dHIS}cm1�P�k_ALM 1O{[� �j4�li0+������r_vb�`  {[��a�R2�nPTCP_VER !{Z�!�_�$EXTL�OG_REQ3v9�i��SIZ����STK���e�~��TOL  m1{Dz;r�A �_BWD�瀠f��R��DI� P�5��Tm1�STEP)�;�nPU��OP_DȌlQF�DR_GRP 19Q{Y�ad 	-�ʟ��P���E%��ڭ?�#���[��� �?
� ������� �!��D�/�h�S��� w��������ѯ
���.��W
$�]�fvM��𜿇�����B�  ��A�  @�3q3��UO���Ϳ��9�$�F�6 F@]�[�g�"σ�~F� ?�  ��ޘ�<P���;O?��9 n���r����q�FEATUROE R�5��Q�ArcTo�ol D�m2E�nglish D�ictionar�yO�4D Sta�ndardH�An�alog I/O�G�AZ�e Shi�ft��rc EQ� Program Select��Softpar�����Weld��ce�dures��@�C�ore��?�Ram�ping��uto���wa'�Upda�teM�matic BackupM��{�ground �EditE�R�Ca�mera��F��C�ell�ܠ�nrR�ndIm���om�mon cali�b UI����sh������c&�.���nYeC�.�ty��s�����n���Moniwtorb�ntr>�eliab��N�D�HCPD۷�ata Acquis��~��iagnosw������ocument Viewe�����ua#�heck Safety	��R�han� Ro-b��rv��qF
�N�ks" F��(�R�xt weavx��chJ�xt. D;IO$�nfiG� wendS Err��QL��s�	r����  �L�FCTN Menu; �  �TP Infa�c(�R�Gen��l�Eq L�]���p Mask EkxcO g�HTJ>��xy Sv#�igh-SpeS �Ski����$�m�municv�on�Hour1�����Mconn}�2�(ncrLstr�uc�M�KAREL Cmd. L��ua�E#Run-;Ti� Env;(�_�+z�sx�S/W�O�License�5"� Book(System)L�MACROs,��/Offse�M�MR����Mec_hStop��t��D���%i���6xS ؔ�x�1>od��wi!t�T8����.$�r;�Optm�?�#��f�il"�'g��%ulti-T�E�P�PCM fun4'��9o��6E�MRe�gi� r��6rib F
KRF��Nu��x��nH��Adju��hN�Ҵ٦MtatupNA�O
Q�RDMU�ot`�scoveLi��Eem0�nw���ERZ� ^ues���9Wo$�_0N�SN�PX b�"H�SNJCli}^��urhӝ_z� %4ujU�o� t1ssag@E�jU�A�{_F� U���!n/IKeMI�LIB;obP F�irm^�%nP1A�cc����TPTX��deln� Xoa�A��%&morIP Simula����fu� P]�j���3�&��ev.eV�r�i3 �oUSB �po���iP� a� bunexcep�tS P(Dbu�uVEC�r��8V���rvo�u�[�{S�PS�C�e
�SUIK�Wx� �8<�b Pl�F X�Z���M��#�FQ�uvn�ԇG�rid
QplayP΍"`��R�r.w���RC�g�100iD/1450���larm Cau�se/Pedj�A�scii��Loa9d" v�Upl����yc��k"Y@Pp@ %�RAp��l�"�NR�TL�oS�Onli?ne Hel���6`L�6L@IA�trG��64MB DRA9M��\�FROe����tl!�0.L�mai�#��[�L%�Sup�mr�1NIР� �cr�o�LS�U��V�Rmi܉�vrt2SK���O�W�i������� ̿ÿտ����%�/� \�S�eϒωϛ��Ͽ� �������!�+�X�O� aߎ߅ߗ��߻����� ����'�T�K�]�� �������������� �#�P�G�Y���}��� ������������ LCU�y��� ����H? Q~u����� ��//D/;/M/z/ q/�/�/�/�/�/�/�/ 	??@?7?I?v?m?? �?�?�?�?�?�?OO <O3OEOrOiO{O�O�O �O�O�O�O__8_/_ A_n_e_w_�_�_�_�_ �_�_�_o4o+o=ojo aoso�o�o�o�o�o�o �o0'9f]o �������� ,�#�5�b�Y�k����� ��Ώŏ׏���(�� 1�^�U�g�������ʟ ��ӟ���$��-�Z� Q�c�������Ư��ϯ �� ��)�V�M�_� ������¿��˿�� ��%�R�I�[ψ�� �Ͼϵ��������� !�N�E�W߄�{ߍߺ� �����������J� A�S��w����� �������F�=�O� |�s������������� B9Kxo ������� >5Gtk}� ����/�/:/ 1/C/p/g/y/�/�/�/ �/�/ ?�/	?6?-??? l?c?u?�?�?�?�?�? �?�?O2O)O;OhO_O qO�O�O�O�O�O�O�O _._%_7_d_[_m_�_ �_�_�_�_�_�_�_*o !o3o`oWoio�o�o�o �o�o�o�o�o&/ \Se����� ���"��+�X�O� a������������ߏ ���'�T�K�]��� ���������۟�� �#�P�G�Y���}��� �����ׯ���� L�C�U���y������� ܿӿ��	��H�?� Q�~�uχϡϫ����� �����D�;�M�z� q߃ߝߧ�������
� ��@�7�I�v�m�� ������������� <�3�E�r�i�{����� ��������8/ Anew���� ���4+=j as������ �/0/'/9/f/]/o/ �/�/�/�/�/�/�/�/ ,?#?5?b?Y?k?�?�? �?�?�?�?�?�?(OO 1O^OUOgO�O�O�O�O��O�O�O�O$_Q � H541�S?Q2DVR782�EW50EUJ614�iW76EUAWSP�QW1�WRCRuX8��VTU�VJ545�iX�VVCAMEUC�LIO�VRI�WU�IFQV6�WCMSyCh�VSTYLiW�2�VCNREQV5�2�VR63PWSC�HEUDOCVqfC�SUEUORS�VR�869iW0tW88�DVEIOfR54�\VR69�VESE�T�W�WJ�YWMG�EUMASKEUPRkXY5h7EVOC�V��`3�X\V�`hXgX5u3�fH^xLCHvwOPLvJ50HvPS�wMC�W�p�g{55tVMDSW�wv;wOP;wMPR�Vpa`0v�`hVPCMg�0��`tW50�5�1�W51P�0�VP�RS�g690vFR=D�VRMCN)f�h�H93hVSNBA�g_wSHLB)fMX߇a`XgNNlx2hVwHTC�VTMI4f�YP�fTPAfTPTX�EL���p�gq8[WYPDVJ95�V�TUT<w950vU�ECvUFR�VV�CC��O�VVIPN4fCSCL��`I�x�tVWEB�VHTT��W6WgWIO��C�G�IG�IPG�S=�RC4fHZXR[66�VR7�gRN�2HvRjz40vu�tV�`DVNVD�fD0���F�CTO�WN�N0vOL'hEND�QVL×SLM�fFVRe XK�]�o��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯��� ������	��-�?�Q� c�u��������� ����)�;�M�_�q� �������������� %7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o	-?Q cu������ ���)�;�M�_�q� ��������ˏݏ�� �%�7�I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ����������'�  �H541)�C�2�H�R782I�50�I�J614y�76^I�AWSPY�1���RCR��8��TU���J545yܘ�V�CAMI�CLIOv�RI�UIFY�=6��CMSCY�گSTYLy�2��C�NREY�52��R�63X�SCHI�DwOCV��CSUI��ORS��R869�y�0��88H�EI�Oh�R54h�R6=9��ESET�۷��J��WMGI�MA{SKI�PRXY��M7I�OC(��3�ܰhڅ�x�w�53�H�LCH��OPLn��J50��PSgcMC��u ��55���MDSW���OP��MPR(�����%�.x�PCMH�0���5051��5u1X0��PRSx��69��FRD�R�MCNy��H93�x�SNBAI�SHLBy�M+����NN(2x�HTC���TMI��e��T{PAh�TPTXi*#EL�u �8g�e��H�J95��TUTv��95��UEC��wUFR�VCC8<�O��VIP��CS�C�*��Ii��WE]B��HTT��6��WIO�:CG�;I�G�;IPGS�:RuC��Hf�R66�ګR7g�RV2��R�&4��5@��U�H�N[VDx�D0�KF�L�CTO��NN��O]Lw�ENDY�LG;wSLMx�FVRh� (�O_a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk }������� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��Ϡ������%�1��STD,�LANGM�H�`�r߄� �ߨߺ��������� &�8�J�\�n���� �����������"�4� F�X�j�|��������� ������0BT fx������ �,>Pbt �������/�/(/:/L/^$RBTL�OPTNu/�/�/8�/�/�+DPNK��/ �/??/?M�$�S?e? w?�?�?�?�?�?�?�? OO+O=OOOaOsO�O �O�O�O�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_�_o#o5o GoYoko}o�o�o�o�o �o�o�o1CU gy������ �	��-�?�Q�c�u� ��������Ϗ��� �)�;�M�_�q����� ����˟ݟ���%� 7�I�[�m�������� ǯٯ����!�3�E� W�i�{�������ÿտ �����/�A�S�e� wωϛϭϿ������� ��+�=�O�a�s߅� �ߩ߻��������� '�9�K�]�o���� �����������#�5� G�Y�k�}��������� ������1CU gy������ �	-?Qcu �������/ /)/;/M/_/q/�/�/ �/�/�/�/�/??%? 7?I?[?m??�?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O��O�O__99�'U�$FEAT_�ADD ?	����TQ\P  	$Xe_w_�_�_ �_�_�_�_�_oo+o =oOoaoso�o�o�o�o �o�o�o'9K ]o������ ���#�5�G�Y�k� }�������ŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;� M�_�q���������˿ ݿ���%�7�I�[� m�ϑϣϵ������� ���!�3�E�W�i�{� �ߟ߱���������� �/�A�S�e�w��� �����������+� =�O�a�s��������� ������'9K ]o���������#5GGTD�EMO RTY   $X�� ������/// &/8/R/\/�/�/�/�/ �/�/�/�/�/+?"?4? N?X?�?|?�?�?�?�? �?�?�?'OO0OJOTO �OxO�O�O�O�O�O�O �O#__,_F_P_}_t_ �_�_�_�_�_�_�_o o(oBoLoyopo�o�o �o�o�o�o�o$ >Hul~��� ����� �:�D� q�h�z�������ݏԏ ��
��6�@�m�d� v�������ٟП�� ��2�<�i�`�r��� ����կ̯ޯ��� .�8�e�\�n������� ѿȿڿ����*�4� a�X�jϗώϠ����� ������&�0�]�T� fߓߊߜ��������� ���"�,�Y�P�b�� ������������� �(�U�L�^������� ���������� $ QHZ�~��� ���� MD V�z����� ��//I/@/R// v/�/�/�/�/�/�/�/ ??E?<?N?{?r?�? �?�?�?�?�?�?
OO AO8OJOwOnO�O�O�O �O�O�O�O__=_4_ F_s_j_|_�_�_�_�_ �_�_oo9o0oBooo foxo�o�o�o�o�o�o �o5,>kbt �������� 1�(�:�g�^�p����� ��ӏʏ܏�� �-�$� 6�c�Z�l�������ϟ Ɵ؟���)� �2�_� V�h�������˯¯ԯ ���%��.�[�R�d� ������ǿ��п��� !��*�W�N�`ύτ� ���Ϻ��������� &�S�J�\߉߀ߒ߿� ����������"�O� F�X��|������ �������K�B�T� ��x������������� G>P}t ������ C:Lyp�� ����	/ //?/ 6/H/u/l/~/�/�/�/ �/�/?�/?;?2?D? q?h?z?�?�?�?�?�? O�?
O7O.O@OmOdO vO�O�O�O�O�O�O�O _3_*_<_i_`_r_�_ �_�_�_�_�_�_o/o &o8oeo\ono�o�o�o �o�o�o�o�o+"4 aXj����� ���'��0�]�T� f������������� ��#��,�Y�P�b��� ������������� �(�U�L�^������� �����ܯ���$� Q�H�Z���~������� �ؿ��� �M�D� Vσ�zόϦϰ����� ���
��I�@�R�� v߈ߢ߬�������� ��E�<�N�{�r�� ������������ A�8�J�w�n������� ��������=4 Fsj|���� ��90Bo fx������ �/5/,/>/k/b/t/ �/�/�/�/�/�/�/? 1?(?:?g?^?p?�?�? �?�?�?�?�? O-O$O 6OcOZOlO�O�O�O�O �O�O�O�O)_ _2___ V_h_�_�_�_�_�_�_ �_�_%oo.o[oRodo ~o�o�o�o�o�o�o�o !*WN`z� �������� &�S�J�\�v������� ���ڏ���"�O�|F�r�  i� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZl~���� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ���������&� 8�J�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x��������������� ,>Pbt� �������(:L^p  qk���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o o&o8oJo\ono�o�o �o�o�o�o�o�o" 4FXj|��� ������0�B� T�f�x���������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ������������ �&�8�J�\�n����� ������������" 4FXj|��� ����0B(Tfvzm� ������/ / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXojo|o�o�o �o�o�o�o�o0 BTfx���� �����,�>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\�n�� ������������� "�4�F�X�j�|����� ����������0 BTfx���� ���,>P bt������ �//(/:/L/^/p/ �/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�?O O 2ODOVOhOzO�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0��B�T�f�x��$FE�AT_DEMOIoN  {������~���INDE�X�������IL�ECOMP S����ޑ�����ԐSETUPo2 Tޕ�?�  N �ѓ�_AP2BCK �1Uޙ  �)y�G�V�%=�z�~��h���{�<�ѯ`� �����+���O�ޯs� �����8�Ϳ߿n�� ��'�9�ȿ]�쿁�� �Ϸ�F���j���ߠ� 5���Y�k��Ϗ�߳� ��T���x����C� ��g��ߋ��,���P� ��������?�Q��� u����(�����^��� ��)��M��q� �6��l� %�2[�� �D�h�/�3/ �W/i/��//�/@/ �/�/v/?�//?A?�/ e?�/�?�?*?�?N?�? �?�?O�?=O�?JOsOt�!�P%� 2:�*.VRzO�O2@*�O�O/C�O_EƮ@PC_H_2@F'R6:3_t^_�_'[T���_�_]U�_�\🐉_o F*.F��OOo1A	_S=o|l8o�o/kSTM�o�o\RbP�o }�o$/kH�oW�gE�0jGIF���e�p��-�0jJPG7��a��eM�
����(ZJS���2@w�ҏ���%
JavaSc�ript�;�CS��h��fU�� %�Cascadin�g Style ?Sheets��@�
ARGNAME�.DTß&L�`\@ן������ğ�DISP*���`�[���*�����H�
T�PEINS.XML˯w�:\߯�����Custom T?oolbar �O��PASSWORD���$NFRS:\�c�"� %Pas�sword Config���?�|� �#�YOG�ֿk�}�� ��0�����f��ϊ�� ����U���y��r߯� >���b���	��-�� Q�c��߇���:�L� ��p������;���_� �����$���H����� ~���7����m�� � ��V�z !�E�i{
� .�Rd��/� /S/�w//�/�/</ �/`/�/?�/+?�/O? �/�/�??�?8?�?�? n?O�?'O9O�?]O�? �O�O"O�OFO�OjO|O _�O5_�O._k_�O�_ _�_�_T_�_x_oo �_Co�_go�_o�o,o �oPo�o�o�o�o? Q�ou��:� ^���)��M�� F������6�ˏݏl� ���%�7�Ə[��� � ���D�ٟh�ҟ� ��3�W�i������ ��ïR��v������ A�Яe���^���*��� N������Ϩ�=�O� ޿s�ϗ�&�8���\� �π���'߶�K���o� ��ߥ�4�����j������#����Y�;��$�FILE_DGB�CK 1U���F���� < �)
SU�MMARY.DG<c��MD:������Diag Summary�����
CONSLO�G������[����Console �log\���	TPOACCNQ���%�������TP Accountin}����FR6:IP�KDMP.ZIP��
'`����E�xception�d��MEMCH�ECK��8�����o�Memory �Data�;�(YF)	FTPN��?�C�q�mment TBDl�;�L =�)ETHERNETa������Ethernet s�?figura���~VDCSVRF`pFXq/�%6 � verify �allt/>�M+=�1%DIFFi/O/�a/�/� %�(d�iff�/�'�6 CHG01�/�/�/{?��!?�?�"*f992 q?X?j?�?
?�?�?@2�3�?�?�?�O �O�O9FVTRNDIAG.LS�OP`OrO_��A ��?nostic_>��T6a)UP?DATES.MP3_~�FRS:\K_��]��Updates List�_��PSRBWLD'.CM�_�wR�_��_p�PS_ROBOOWEL����AHADOW�O�O�O��o�Shado�w Change�s�oqQbNOTI;/lo~o��Notificx"�o;�+@AG�� j�9����� w���B��f�x� ���+���ҏa����� ���'�P�ߏt���� ��9�Ο]�����(� ��L�^�ퟂ����5� ��ܯk� ���$�6�ů Z��~������C�ؿ �y�ϝ�2���?�h� ����ϰ���Q���u� 
�߫�@���d�v�� ��)߾�M����߃�� ��<�N���r���� 7���[������&��� J���W������3��� ��i�����"4��X ��|��A�e ��0�Tf� ���O�s/ /�>/�b/�o/�/ '/�/K/�/�/�/?�/ :?L?�/p?�/�?�?5? �?Y?�?}?�?$O�?HO �?lO~OO�O1O�O�O gO�O�O _2_�OV_�O z_	_�_�_?_�_c_�_ 
o�_.o�_Rodo�_�o o�o�oMo�oqo�o <�o`�o��% �I����8� J��n����!���ȏ W��{��"���F�Տ j�|����/�ğ֟e� �������+�T��x� �����=�үa���� ��,���P�b�񯆿� ��9����o�ϓ�(� :�ɿ^��ϔ�#ϸ� G�����}�ߡ�6����C�l�N��$FIL�E_FRSPRT�  ��V�������M�DONLY 1U���N� 
 ��)MD:_VD�AEXTP.ZZ�Zs�$���
�6�%NO Back file ��N�S�6�\��� ��Iߍ������i��� ���4���X�j���� �����S���w��� B��f����+ �O����> P�t�'�� ]��/(/�L/� p/�//�/5/�/�/��?VISBCK�؝�>��*.VD�/'?�� FR:\� I�ON\DATA\�?�"� Vis?ion VD(�S? a/�?�?�/�?�/�?�? O+O�?OO�?sO�OO �O8O�O\OnO_�O'_ 9_�O]_�O�__�_�_ F_�_j_�_o�_5o�_ Yo�_�_�oo�o�o�o �oxo�oC�og �o��,�P�t���{�LUI_C�ONFIG V��	1&� $ ���q��������ˏݏ��$ |x ��!�3�E�W�g��� ��������ҟi��� �,�>�P��t����� ����ίe����(� :�L��p��������� ʿa�� ��$�6�H� ߿l�~ϐϢϴ���]� ����� �2�D���h� zߌߞ߰���Y����� 
��.���?�d�v�� ���C��������� *���N�`�r������� ?�������&�� J\n���;� ���"�FX j|��7��� �//�B/T/f/x/ �/!/�/�/�/�/�/? �/,?>?P?b?t?�?? �?�?�?�?�?O�?(O :OLO^OpO�OO�O�O �O�O�O _�O$_6_H_ Z_l_~__�_�_�_�_ �_�_�_ o2oDoVoho zoo�o�o�o�o�o}o �o.@Rd�o� �����y�� *�<�N�`�������� ��̏ޏu���&�8� J�\�󏀟������ȟ ڟq����"�4�F�X� �|�������į֯f���|�$FLU�I_DATA �W�����j���RES�ULT 2X��0� �T�� �L�^�p��������� ʿܿ� ��$�j�9� L�^�pςϔϦϸ��π���� ��$�6�G�?�j�0���~�i�{��r��߱� ����������/�A� S�e�w�6Îߡ���� ��������1�C�U�g�y�j�
�yߟ�]� ��������
.@ Rdv����� ���*<N` r�������� ��/��8/J/\/n/�/ �/�/�/�/�/�/�/? "?�F?X?j?|?�?�? �?�?�?�?�?OO� ?O/cO%/'O�O�O�O �O�O�O__,_>_P_ b_t_3?�_�_�_�_�_ �_oo(o:oLo^opo /O�oSO�o�o�_�o  $6HZl~� ����_��� � 2�D�V�h�z������� �o�o�o���o@� R�d�v���������П ������<�N�`� r���������̯ޯ� ��ӏ���A�k�-� ������ȿڿ���� "�4�F�X�j�)��Ϡ� ������������0� B�T�f�%�7�I�[��� �������,�>�P� b�t�����{��� ����(�:�L�^�p� �����������ߛ߭� ��6HZl~� �������� 2DVhz��� ����
//���� ��a/#�/�/�/�/�/ �/�/??*?<?N?`? q?�?�?�?�?�?�? OO&O8OJO\OnO-/ �OQ/�Ou/�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�O�_�_oo0o BoTofoxo�o�o�o�o O�o�O�O,>P bt������ ����_:�L�^�p� ��������ʏ܏� � ��o3��oW���� ����Ɵ؟���� � 2�D�V�h�'������� ¯ԯ���
��.�@� R�d�#���G������ �����*�<�N�`� rτϖϨϺ�y����� ��&�8�J�\�n߀� �ߤ߶�u�������� Ͽ4�F�X�j�|��� �������������0� B�T�f�x��������� �����������5 _!������ �(:L^� ������� / /$/6/H/Z/+= O�/s�/�/�/? ? 2?D?V?h?z?�?�?�? o�?�?�?
OO.O@O ROdOvO�O�O�O�O}/ �/�/_�/*_<_N_`_ r_�_�_�_�_�_�_�_ o�?&o8oJo\ono�o �o�o�o�o�o�o�o �O�O�OU_|�� �������0� B�T�oe��������� ҏ�����,�>�P� b�!��E��iΟ�� ���(�:�L�^�p� ��������ɟܯ� � �$�6�H�Z�l�~��� ����s�տ������ � 2�D�V�h�zόϞϰ� ��������
�ɯ.�@� R�d�v߈ߚ߬߾��� �����ſ'��K�� ����������� ��&�8�J�\�߀� �������������� "4FX�y;� �s����0 BTfx���m� ���//,/>/P/ b/t/�/�/�/i�� �/?�(?:?L?^?p? �?�?�?�?�?�?�? O �$O6OHOZOlO~O�O �O�O�O�O�O�O�/? �/)_S_?z_�_�_�_ �_�_�_�_
oo.o@o RoOvo�o�o�o�o�o �o�o*<N_ _1_C_�g_��� ��&�8�J�\�n��� ����coȏڏ���� "�4�F�X�j�|����� ��q������0� B�T�f�x��������� ү������,�>�P� b�t���������ο� ��ß՟�I��p� �ϔϦϸ������� � �$�6�H��Y�~ߐ� �ߴ���������� � 2�D�V��w�9ϛ�]� ��������
��.�@� R�d�v����������� ����*<N` r���g����� ��&8J\n� ��������� "/4/F/X/j/|/�/�/ �/�/�/�/�/�?� ???x?�?�?�?�? �?�?�?OO,O>OPO /tO�O�O�O�O�O�O �O__(_:_L_?m_ /?�_�_gO�_�_�_ o o$o6oHoZolo~o�o �oaO�o�o�o�o  2DVhz��]_ �_�_���_�.�@� R�d�v���������Џ ��o�*�<�N�`� r���������̟ޟ� ����G�	�n��� ������ȯگ���� "�4�F��j�|����� ��Ŀֿ�����0� B���%�7���[��� ��������,�>�P� b�t߆ߘ�W������� ����(�:�L�^�p� ����e�wω���� �$�6�H�Z�l�~��� ������������  2DVhz��� ����������= ��dv����� ��//*/</��M/ r/�/�/�/�/�/�/�/ ??&?8?J?	k?- �?Q�?�?�?�?�?O "O4OFOXOjO|O�O�O �?�O�O�O�O__0_ B_T_f_x_�_�_[?�_ ?�_�?oo,o>oPo boto�o�o�o�o�o�o �o�O(:L^p ��������_ ��_3��_�l�~��� ����Ə؏���� � 2�D�h�z������� ԟ���
��.�@� �a�#�����[���Я �����*�<�N�`� r�����U���̿޿� ��&�8�J�\�nπ� ��Q���u����ϫ�� "�4�F�X�j�|ߎߠ� �������ߧ���0� B�T�f�x������ ����������;��� b�t������������� ��(:��^p �������  $6����+�� O������/ / 2/D/V/h/z/�/K�/ �/�/�/�/
??.?@? R?d?v?�?�?Yk} �?�OO*O<ONO`O rO�O�O�O�O�O�O�/ __&_8_J_\_n_�_ �_�_�_�_�_�_�?�? �?1o�?Xojo|o�o�o �o�o�o�o�o0 �OAfx���� �����,�>��_ _�!o��Eo����Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� O���s�կ����� � 2�D�V�h�z������� ¿Կ濥�
��.�@� R�d�vψϚϬϾ��� �ϡ��ů'����`� r߄ߖߨߺ������� ��&�8���\�n�� ������������� "�4���U��y���O� ����������0 BTfx�I�� ���,>P bt�E���i��� ��//(/:/L/^/p/ �/�/�/�/�/�/� ? ?$?6?H?Z?l?~?�? �?�?�?�?���O /O�VOhOzO�O�O�O �O�O�O�O
__._�/ R_d_v_�_�_�_�_�_ �_�_oo*o�?�?O O�oCO�o�o�o�o�o &8J\n� ?_������� "�4�F�X�j�|���Mo _oqoӏ�o����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ����Ï%��L�^�p� ��������ʿܿ� � �$��5�Z�l�~ϐ� �ϴ���������� � 2��S��w�9��߰� ��������
��.�@� R�d�v��߬���� ������*�<�N�`� r���Cߥ�g������� &8J\n� �������� "4FXj|�� ��������/�� �T/f/x/�/�/�/�/ �/�/�/??,?�P? b?t?�?�?�?�?�?�? �?OO(O�IO/mO OC?�O�O�O�O�O _ _$_6_H_Z_l_~_=? �_�_�_�_�_�_o o 2oDoVohozo9O�O]O �o�o�O�o
.@ Rdv����� �_���*�<�N�`� r���������̏�o�o �o��#��oJ�\�n��� ������ȟڟ���� "��F�X�j�|����� ��į֯�����ݏ ���u�7������� ҿ�����,�>�P� b�t�3��Ϫϼ����� ����(�:�L�^�p� ��A�S�e��߉��� � �$�6�H�Z�l�~�� ����������� � 2�D�V�h�z������� �����ߥ߷���@ Rdv����� ����)N` r������� //&/��G/	k/- �/�/�/�/�/�/�/? "?4?F?X?j?|?�/�? �?�?�?�?�?OO0O BOTOfOxO7/�O[/�O /�O�O__,_>_P_ b_t_�_�_�_�_�_�? �_oo(o:oLo^opo �o�o�o�o�o�O�o�O �O�oHZl~� ������� � �_D�V�h�z������� ԏ���
���o=� �oa�s�7�������П �����*�<�N�`� r�1�������̯ޯ� ��&�8�J�\�n�-� w�Q���ſ������ "�4�F�X�j�|ώϠ� ���σ�������0� B�T�f�xߊߜ߮��� �ɿ�����ٿ>�P� b�t��������� ������:�L�^�p� ��������������  �������i+� ������  2DVh'���� ����
//./@/ R/d/v/5GY�/} �/�/??*?<?N?`? r?�?�?�?�?y�?�? OO&O8OJO\OnO�O �O�O�O�O�/�/�/_ �/4_F_X_j_|_�_�_ �_�_�_�_�_o�?o BoTofoxo�o�o�o�o �o�o�o�O;�O _!_������ ���(�:�L�^�p� �������ʏ܏� � �$�6�H�Z�l�+�� O��s؟���� � 2�D�V�h�z������� ¯�����
��.�@� R�d�v���������}� ߿���şǿ<�N�`� rτϖϨϺ������� ��ӯ8�J�\�n߀� �ߤ߶���������� Ͽ1��U�g�+ߎ�� ������������0� B�T�f�%ߊ������� ������,>P b!�k�E��{�� �(:L^p ����w��� / /$/6/H/Z/l/~/�/ �/�/s���/?� 2?D?V?h?z?�?�?�? �?�?�?�?
O�.O@O ROdOvO�O�O�O�O�O �O�O_�/�/�/�/]_ ?�_�_�_�_�_�_�_ oo&o8oJo\oO�o �o�o�o�o�o�o�o "4FXj)_;_M_ �q_�����0� B�T�f�x�������mo ҏ�����,�>�P� b�t���������{� ���(�:�L�^�p� ��������ʯܯ� � ���6�H�Z�l�~��� ����ƿؿ����͟ /��S��zόϞϰ� ��������
��.�@� R�d�uψߚ߬߾��� ������*�<�N�`� ρ�Cϥ�g������� ��&�8�J�\�n��� ������u������� "4FXj|�� �q�������0 BTfx���� ���/��,/>/P/ b/t/�/�/�/�/�/�/ �/?�%?�I?[?/ �?�?�?�?�?�?�? O O$O6OHOZO/~O�O �O�O�O�O�O�O_ _ 2_D_V_?_?9?�_�_ o?�_�_�_
oo.o@o Rodovo�o�o�okO�o �o�o*<N` r���g_�_�_� ��_&�8�J�\�n��� ������ȏڏ����o "�4�F�X�j�|����� ��ğ֟������ �Q��x��������� ү�����,�>�P� �t���������ο� ���(�:�L�^�� /�A���e������� � �$�6�H�Z�l�~ߐ� ��a���������� � 2�D�V�h�z���� oρϓ�����.�@� R�d�v����������� ������*<N` r������� ��#��G	�n� �������/ "/4/F/X/i|/�/�/ �/�/�/�/�/??0? B?T?u?7�?[�? �?�?�?OO,O>OPO bOtO�O�O�Oi/�O�O �O__(_:_L_^_p_ �_�_�_e?�_�?�_�? �_$o6oHoZolo~o�o �o�o�o�o�o�o�O  2DVhz��� �����_��_=� O�v���������Џ ����*�<�N� r���������̟ޟ� ��&�8�J�	�S�-� w���c�ȯگ���� "�4�F�X�j�|����� _�Ŀֿ�����0� B�T�f�xϊϜ�[��� ����ϵ��,�>�P� b�t߆ߘߪ߼����� �߱��(�:�L�^�p� ������������ ������E��l�~��� ������������  2D�hz��� ����
.@ R�#�5��Y��� ��//*/</N/`/ r/�/�/U�/�/�/�/ ??&?8?J?\?n?�? �?�?cu��?�O "O4OFOXOjO|O�O�O �O�O�O�O�/�O_0_ B_T_f_x_�_�_�_�_ �_�_�_�?o�?;o�? boto�o�o�o�o�o�o �o(:L]op ������� � �$�6�H�oi�+o�� Oo��Ə؏���� � 2�D�V�h�z�����] ԟ���
��.�@� R�d�v�����Y���}� ߯�����*�<�N�`� r���������̿޿� ���&�8�J�\�nπ� �Ϥ϶������ϫ�� ϯ1�C��j�|ߎߠ� ������������0� B��f�x������ ��������,�>��� G�!�k���W߼����� ��(:L^p ��S����  $6HZl~� O���s�����/ / 2/D/V/h/z/�/�/�/ �/�/�/�
??.?@? R?d?v?�?�?�?�?�? �?����9O�`O rO�O�O�O�O�O�O�O __&_8_�/\_n_�_ �_�_�_�_�_�_�_o "o4oFoOO)O�oMO �o�o�o�o�o0 BTfx�I_�� �����,�>�P� b�t�����Woio{oݏ �o��(�:�L�^�p� ��������ʟܟ�� �$�6�H�Z�l�~��� ����Ưدꯩ��͏ /��V�h�z������� ¿Կ���
��.�@� Q�d�vψϚϬϾ��� ������*�<���]� ���C��ߺ������� ��&�8�J�\�n�� ��Q϶���������� "�4�F�X�j�|���M� ��q����ߗ�0 BTfx���� ����,>P bt������ ��/��%/7/�^/p/ �/�/�/�/�/�/�/ ? ?$?6?�Z?l?~?�? �?�?�?�?�?�?O O 2O�;//_O�OK/�O �O�O�O�O
__._@_ R_d_v_�_G?�_�_�_ �_�_oo*o<oNo`o ro�oCO�OgO�o�o�O &8J\n� ������_�� "�4�F�X�j�|����� ��ď֏�o�o�o�o-� �oT�f�x��������� ҟ�����,��P� b�t���������ί� ���(�:����� �A�����ʿܿ� � �$�6�H�Z�l�~�=� �ϴ���������� � 2�D�V�h�zߌ�K�]� o��ߓ���
��.�@� R�d�v������� ������*�<�N�`� r��������������� ����#��J\n� ������� "4EXj|�� �����//0/ ��Q/u/7�/�/�/ �/�/�/??,?>?P? b?t?�?E�?�?�?�? �?OO(O:OLO^OpO �OA/�Oe/�O�/�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�?�_o o 2oDoVohozo�o�o�o �o�o�O�o�O+�_ Rdv����� ����*��_N�`� r���������̏ޏ�� ��&��o/	S�}� ?����ȟڟ���� "�4�F�X�j�|�;��� ��į֯�����0� B�T�f�x�7���[��� Ͽ������,�>�P� b�tφϘϪϼ��ύ� ����(�:�L�^�p� �ߔߦ߸��߉����� ��!��H�Z�l�~�� ������������ � ��D�V�h�z������� ��������
.�� ���s5���� ��*<N` r1������� //&/8/J/\/n/�/ ?Qc�/��/�/? "?4?F?X?j?|?�?�? �?�?��?�?OO0O BOTOfOxO�O�O�O�O��O�/�O�/_%Y�$�FMR2_GRP� 1Y%U�� �C4 w B��0	 �0�c_u\`PF�6 F@�S�Q�T�J`Sx�_�]`P?�  �_��_<P�a;O?��9 n�e�]�A`+o=kBH]SB�YPX`;a@�33�ce�\�_�o�Y@UO߯a�o�_�o�o�o �o4XC|g����}9R_CF�G ZF[T ���(�:��{NO� FZ
F0�p� u��|RM_C�HKTYP  �6Q�0NPPPP8QRO=M��_MIN���3W�����|`X9P�SSB�s[%U aV��5��
���uTP_D�EF_OW  ��4NS1�IRCO�M��B��$GENOVRD_DO����1o�THR�� �d��du�_ENB�a� u�RAVC�?S\Ӈހ �@�U"���1��?��P�sj �ՑOU*BPbF\x�sXF�nsU<�� �]�ǯq������3C�
YP�YP�%��d��1A@M�?�U�vY��\#�֐SMT?Sc��RP��4��$HOS�TC�r1dFY߀[��? 	
�
˓
��6:��9eVχϙϫϽ���uπ�� ��$�G�H���	�anonymou�sK�yߋߝ߯���  	��-�
�A�c���R� d�v���Ϭ������ ���M�_�<�N�`�r� ������������7� &8J\��� �����!�3�" 4FX�������� ���//e// T/f/x/�/��/��/ �/�/??as�� �/s?��?�?�?�?�? 9/O(O:OLO^O�?�/ �/�O�O�O�O�O5?G? Y?_mOZ_�?~_�_�_ �_�_q_�_�_o oC_ Do�Ohozo�o�o�o�O 	__-_
Aoc_@R dv��_���� �Mo_o<�N�`�r� ���o�o�o���7 �&�8�J�\������ ����ُǟ!����"��4�F����ENT {1e�� P!ڟ.��  ����ï ��篪��ί/��;� �d���L���p�ѿ�� �����ܿ�O��s� 6ϗ�Zϻ�~ϐ��ϴ� ���9���]� �Vߓ� �߷�z��ߞ������ ��4�Y��}�@��d� ����������C���g�*�QUIC�C0t�P�b�����1 ��������2���c!ROUT�ERd@R�!�PCJOG���!192.16?8.0.10����?CAMPRT��!�1� +R�T}/A�h�NA�ME !u�!�ROBO�S_�CFG 1du�� �Au�to-start{ed��FTP��;!͏ϟf/��/�/ �/�/�/o��/??,? O/=?�/t?�?�?�?�? ��/&/8/OL?n/,O ]OoO�O�OZ?�O�O�O �O�O"O�O5_G_Y_k_ }_�_������ʏ_�_ BOo1oCoUogo._�o �o�o�o�o�_xo	 -?Qc�_�_�_� �o�o���)��o M�_�q������:��� ݏ���%�l~� ��������ǟٟ� ��ď!�3�E�W�i��� �����ïկ���@� R�d�A�x�e������� ������|�����+� N�O��sυϗϩϻ� ��&�8�:��n�K� ]�o߁ߓ�ZϷ����� ����"ߤ�5�G�Y�k� }�������Ϩ���� B��1�C�U�g�.�� ����������x�	�-?Q��_ER�R f�aqP�DUSIZ  j��^���>�?WRD ?%����  guest�����);�SCD_�GROUP 3g�, !��] �LOA���RES�TM�� $�T_�EN�Bs TTP_AU�TH 1h� �<!iPendCanGR.���A�!KAREL:q*R/[/m-KC�/��/�/z VISI?ON SETk?�/F!??1?w#U? C?m?g?�?�?�?�?�?��>!$CTRL �i�;H��
��FFF9E3�?���FRS:DE�FAULT`L�FANUC We�b Server `JNB!$��	L�O�O��O__,_oWR_�CONFIG ]jp�`O�qIDL_CPU�_PC@��B�����P BH�UMI�N�\x�UGNR_�IOz�����PN�PT_SIM_D�O�V�[STAL�_SCRN�V ��6F�QTPMODN�TOLg�[�ARTY�X�Q�V� %  g�x�SOLNK 1k�}�o�o�o��o�o �bMAS�TE�Pzi�UOSLAVE l��AuRAMCACH�E0(bO'!O_CcFGr�c�sUO0<��rCYCLq�u�y@_ASG 1maW�
 �)� ;�M�_�q����������ˏݏ��{�rNU�M��	
�rIP�o�wRTRY_C�N@�R�
�ra_USPD��a�� �r�p�rnP~u��u��PSDT_ISO_LC  P{v"~�J23_DSrd�.N�OGg1onP{<��d<�P�� ?��R��?��館Q��̯ޯ�@���&�8�J�����@��*��P�qi��Php�ECso�UKANJ�I_*pK�_³� MON pp;_��y�(�:�L�^�pϒ$~"��qa\EF�ŭ���CL_L�P'�J��İEYLOGGI�N�pu�F����$LANGUA�GE �Fab�yD <�qLG�qyr�y�a ���xu �e����P�V��'0�����;���cMCH ;��
���(UT1:\���� �������� �!�3�E�\�i�{���(���lLN_D?ISP sP�ؘ������OC4b�RD�z�S�A@�OGB�OOK tM�d`��>A���k�X�� ����������<O�Y���	>F	Q����Й�N`��O�_B�UFF 1u�me2kE�j�FB� iG��G> P}t�������///C/��~D�CS w�{�=���G��/�/�/�/Z$IO 1x�{ ğ3D��?*?<?N?b?r?�? �?�?�?�?�?�?OO &O:OJO\OnO�O�O�Oh�O�O�%E�PTM�dh�#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o-�N�BSEV�����FTYP�_�o�m��RSh���|>��FL 2y=����/�������(TP����b}'�NGNAM��6%.�V$UPS��G�Ih�����f�_L�OADPROG �%��%REQ�MENU��MA?XUALRM'��A85�̀l�_PRh���� E�	ˀC��z�M�������,�P �2{� ت	Z�aڀ	�|�f4� �~����������(Ο ���3��(�i�T��� x���ï���ү��  �A�,�e�P�����~� �����ƿؿ��=� (�a�s�VϗςϻϞ� ������� �9�K�.� o�Zߓ�v߈��ߴ��� ���#��G�2�k�N� `������������ �
�C�&�8�y�d��� ������������ć�DBGDEF �|$�:!"�$6 _L?DXDISAQ�#���#MEMO_AP�K�E ?$�
 H�������"ˀISCW 1}$�%�� oy�M�����QE_MSTR �~�m%SCD 1���T/�x/ c/�/�/�/�/�/�/�/ ??>?)?b?M?r?�? �?�?�?�?�?O�?(O O%O^OIO�OmO�O�O �O�O�O _�O$__H_ 3_l_W_�_{_�_�_�_ �_�_o�_2ooBoho So�owo�o�o�o�o�o �o�o.R=va ����������<�'�`��MJPTCFG 1�+�]�%�����MI/R 1�%Ԁp�@T�q���T��< G ?� �%��t�7�q�� i������������� 1�C�֟��j�L�V�x� ��P�����ί��0� T�E �q����8��� ������򿐿����  �B�p�R��ϵ���Z� |���п����6���>� l�R�d߆߈ߖ����� �ߞ���2���@�z� `����������� +�=��������X�b� t�������������* ��o�6��� ������
 @nP���Xz ����4/�,/j/@P/b/�/�/���K��;���  �/���LTARM_�"�̅� �"����6?�>4��METPU ; T����%���NDSP_ADC�OLX5� c>CMN�Ty? l5MST ��-�?���!�?|�4l5POSCF�7=�>PRPM�?�9[STw01���4܁<#�
gA[�gEwO �GcO�O�O�O�O�O�O _�O_G_)_;_}___�q_�_�_�_�_�Ql1S�ING_CHK � |?$MODAQ3����,�.#e�DEV 	��	�MC:WlHSI�ZEX0�-�#eTA�SK %��%$�12345678�9 �o�e!gTRI������ l̅% &�O2}���c�YP�a��9d"cE�M_INF 1��7;a`)AT&FV0E0X��})�qE0V1�&A3&B1&D�2&S0&C1S�0=�})ATZ�#�
�H'�O��qCw��A���b�ˏ���� �&���� ���3���ۏȟڟ�� ����"�4��X��� ��A�S�e�֯៛�� C�0����f�!���q� ����s�俗�����ͯ >��bϙ�sϘ�K��� w��������ɿۿL� ���#ϔߦ�Y���� �ߩ߳�$���H�/�l� ~�1ߢ�U�g�yߋ��� �� �2�i�V�	�z�5����������PoNIT�OR�0G ?kk �  	EXESC1�223E45�`789�� �(�4�@� L�X�d�p�T|�2�2�2�U2�2�2�2�U2�2�2�3��3�3(#aR_G�RP_SV 1��{ (�Q���#aƮa_Ds�n�IO/N_DB-`�1m�1  ��0dKc"%p0&��2Gg���N Bl"%"Fi-ud1}e�/�/�/1�PL_NAME �!�e� �!�Default �Personal�ity (fro�m FD)b"P0R�R2� 1�L?68L@P�!K`
 d�:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O�O�Oc(2)?�O�O�O __,_>_P_b_t_f"<�O�_�_�_�_�_�_ 
oo.o@oRodotl�"�Q �_�m
�o�of$P �o�o $6HZ l~������ ��o�o2�D�V�h�z� ������ԏ���
� �.�@��!�v����� ����П�����*�@<�N�`�r�����e�����ïխf"d����(�6�������y�d���P� ������Ŀֿ������:ϐ��]�m�f"��	`���ϲ��σ�:�oAb)������c' A� � /�	23��)X ����E ���X, �@D�  t�?��z�n�?f |�f!AI��t�j��;�	�l��	 �� � �h�Y Z ����� � x � �� ��Ґ�K_�K }K7X��K��J��?J�+Ƀ�%���ԯC@�6@��
�\��(E@��Sє��.��=�N��������T;f�a������$��* � ´  �@ �>�����z�w�����<�
�����Z!�/�����yD� � �  � W �`�#  �l�����-�	'� �� ��I� ��  �0�&�:��È��È=�s����x�@��@��%�f���f�(��2�+�a!v  '��Y��@!�p@����@��@��@���C��C� �W� C��C��C��R!�A��������%"T�Bb $/�0�Lf!Dz��o ��~������R!���A �кD� � X ,f �?��ffG�*/</� }�q/�+�8~`�/�*�>��$��(�(~`�%P�(�������>�$��ܴ<��	<S�;��9<��<#*�o<��M,@�K;|��f��",��?fff? ?&��0T�@�.�2�?J<?N\��55	 ��1��(�|��?z��? j7��[/0OOTO?OxO cO�O�O�O�O�O�O{h�5F���O2_�OV_ �?w_�9I_�_E_�_�_ �_�_oooLo7opo [o�oo�o�oU�o�o ��m_3�_Z�o~���O*��& Q/�wl��q
�m.��+�d�V���Aa0��5u�CP���L�č?Ƀ���#��Yĭ/Ӄ6�B]�D���CC3� z����ؼ����@I�l�����A��A���PA �R?��1>�-8������ÍO\������Q���#�
؞����AиRA����C;����Q섟"\)�C0���q�Bo
=��Q�����8�Hp���G� H�0��H��E1�� C�&�Hy���I��H��%F�� E,�s��]�i�EI��@�H���H��E# D�7� د�կ���2��V� A�z�e�w�����Կ�� �����@�R�=�v� aϚυϾϩ������� ��<�'�`�K߄�o� �ߺߥ��������&� �J�5�G��k��� ��������"��F� 1�j�U���y������� ������0T? x�u�����@�P�(<g3�(��	4���<�̷�t�Ӂ�3�� ����ʭ��Ӂ� &�n�
/4�f4yϱ$-$)d/R/�/Pv/�/�,ՅPD2P�.�a�o?Z?=?(?a?L<?g?n?�?�?�?��?�?  ���� �?�?+OOOO:OsO? �o�O�O�O�L7�O�O�_�O _F_4_JQ� L_^_�_�_�_�_�_�Z�  2jOo  B(��}���Cq���Ӏ@��Rodovo�o�o�o�mۃo�o�o�/AӄhDӀ�Ӏ�aӀ؎
 I������ ��)�;�M�_�q�����sq ���1���"�$MSKCFMAP  $%� �V�sqoq莼�ONREoL  �%Ӂ��P��EXCFEN�B�
у���FN�y�'��JOGOV�LIM�d��d���KEY�q�z�_PAN��������RUNa���S?FSPDTY� '�<���SIGN���T1MOTc�����_CE_GRP� 1�$%Ӄ\ dOh�\O�����T��ɯ �����#�گG��� <�}�4�����j�׿�� ���Ŀ1��*�g�� �ϝτ���x����������f��QZ_ED�IT�͇��TCO�M_CFG 1�Bɍ~vv߈ߚ�
V�__ARC_"��%�P�T_MN_MO�DE��0�UA�P_CPL��4�N�OCHECK ?=ɋ �%� 3�E�W�i�{���� ����������/�A���NO_WAITc_L�K�6�NT^���ɋu|��_ER�R@�2�ɉ�Q� A��������X4F��MO�����|ߍ�5<���?����np���_PARAM��ɋ�rv�3u7�_�^ =�P345678901x�� s����//�09/K/'+t7�}/�,�"�/��ODRDS�P���0�OFFS?ET_CARA����&DIS�/�#S_�A��ARK�L�O�PEN_FILE�0h���Lִ�OPT?ION_IO�����m0M_PRG %Ɋ%$*�?�>I3�WO50�F�B0� �5���2���0@�'A	 ����C���#�� R�G_DSBL  �Ʌ�v|rO�!R�IENTTO���!C�mpҁ,a� UT_SIM_Du7�Ђ��� V� LCT ���H��4����I�%y��A_PEX���?TRAT�� �d0�T� UP S��N�pK��i_ {_XrfS`�gq�Rn��}]�$�2?��L68L@P�C
 d�/�_o o*o<oNo`oro�o�o �o�o�o�o�o&8J\��2�_�� �����
��.� �{X�j�|������� ď֏�������� �G�X��PX�~��"P k�����̟ޟ��� &�8�J�\�n������� ����������"�4� F�X�j�|�������Ŀ ֿ���ɯۯ0�B�T� f�xϊϜϮ������� ����,�>���|C�}ߏ�S�$�� �ޤ�����b�bݢ/3��W�
�@L�v�l� ~��������J��Q0�'�)L�	``�Z�xl�~���:�o�A���������K�A��  ���T�POOP1��[�v���TH��E�=DX,? @D�  2�4�,?�D442�9�h;�	l�	�@� � �h�� ��� � x? � � ��J��H�H2�-�HL��H�l�H�WG����=�3Ho��J�C�R�@p�@ז@�PT1w#��0@�S �>PP%ICUB��<��K�`�@��a�y��  �  _�  � #�0��*&�H/�	'�� � f"I� �  ����=��͊/�+�@�/� �>A�/DM+>B���N�@4?  'x0L4�0}C�@C�� C�C�C�Y?k?D� � �A�!�������/��B�@�1 �����!
ENz�-O �QO<OaO�O^/p(�1<�E�S� �<��1��P.   �?�faf��O�O�O 7��/_A[sA8�W_eZ>��' �FjJ(��UP�X�I�����#�T[ܾ<��	<S�;��9<��<#*�o<��5�\@�	k:��#�R���?fff?� ?&�D`oD@�.Vb�?J<?N\�be:� �2?aKjI:�o8�o (g~_�o�o�o6 !ZE~�{�� �����o�o�o� h����w�����ԏ�� я
���.��R�=�v� a�?��o�e+��O�����<�N�`�r�Z���@_��l� /�ȯ�+��ׯ�"����A`>��?�C�s�
�<П��?�ء�����̿n	�/X�j��B�D90CC��ޚ�������^�@I��*����A���A��PA ��R?�1>��-���������O\����Q����#�
�����A�иRA���C;���Q�B���0\)C0����qBo
=���Q�������Hp��G�� H�0�H��E1� C����Hy��I���H��%F�� �E,�1߯i�E�I��@H����H��E# D����ߨߓ��� ���������8�#�5� n�Y��}������� �����4��X�C�|� g��������������� 	B-fxc� ������ >)bM�q�� ���/�(//L/ 7/p/[/m/�/�/�/�/ �/�/?�/6?H?3?l? W?�?{?�?�?�?�?�?tO��(��3�([���T��BE�5�̷�2ODOX�3���8^OpO~B�ʭ�O�O�X�� &n�O�O4�f4yϱ�M �I"__F_4_j_X\��%PbP�^�����_@O�_�_�_o
l?%o�,oeoPouo�o�o  ���ʞo�o�o�o �o1�_��dR�v|7����������
��R�@�pv�d�����  2(�я  BG�;�G�C/�D�X�@K��"�@4�F�X�j�{����������ɟ۟���X�J��X�X���X���
 �W�i� {�������ïկ������/�A���1� ����K1��"�$�PARAM_ME�NU ?�E��  �MNUTOOL�NUM[1]݆���F~������AWEPCR��.�$INCH_RA�TE��SHEL�L_CFG.$J�OB_BAS߰ �WVWPR.�$CENTER_�RI������AZI�MUTH OPT�B����ELEV�ATION TCگ���DW�TY�PE SN�AR�CLINK_AT~ �STATUSǳ~]�__VALU߱�̰LEP��.$WP_�����U�̢� �����������7�2��D�V��z�SSREL_ID  �E��Q���USE_P�ROG %��%x{��ߏ�CCRT����Q����_HOST7 !��!��5���T�P��Q��*��S����_TIMEsOU�Ս�  z�?GDEBUG�Љ����GINP_FLgMSK����TR����PGd�  ����$�CH����Q���z�tߪ����� ����(:c^ p�������  ;6HZ�~ ������//� /2/[/��WORD� ?	��
 	�RS�CPN<n�BMAIW��#3SU&��#TEt�C�STYL C�OL0eW(�/W�TR�ACECTL 1��E�� ��P�P7DT Q��ED0!0D �� �S��QQ6�[;q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#��5�G�Y�k�}�6LE�W���5��3  ��6_UP ��<;b������ ���&�0�M$a���R�\0R�  ���)_DEFSPD� ���2�� � �z�INؐT�RL ���a�8�!�h�PE_CON�FIܐ�7�t��M!b,LIDٓ����	ĨGRP �1�9 l�M!A>ff���\�
=D�  DZ� D
�-@�
�M d!�?�O�������H�"�$�i� ´����m�B��̱�������̿���&�B34�$�]�o�Y� <<j��tϭ�pϪ��� ����ό��O��_߈��p��z�ӳ�M 
 ���ߊ������5� � Y�D�}�h�������������*�)<��
V7.10be�ta1�� A��k�\�B
��(�Y�?&ffp�>�.{X�
���{��X�B!념�?A{33A�&�(�h� -�����������pM"��3E�WM$ғ�KNOW_M  0��Ȥ�SV �:�%��������IM"G��M��=�(�	�����.�*~ ����M#�)�Y�@)���`M % .ѐȡMR��=�$����f/x+���ST�1 1�<9^ 4�()� o��/�/�/
?�/?!? S?E?W?�?{?�?�?�? �?O�?�?>OO/OtOSOeOwO�'2�,��/����<�O�O� 3 �O�O�O�O�'4_-_?_Q_�'5n_�_�_�_��'6�_�_�_�_�'7 o&o8oJo�'8goyo��o�o�'MAD�� �ȕ�EOVLD � ���P}�$P�ARNUM  p�+?Q�#SCHy ȕ
�wlq�y��uUPDl=u��>�E_CMP_u�����_�'ݥ%�ER/_CHK3�ۣ �G�0�B�RSA �ȡG_MOp����_��~�E_RES_G� ���
��p�"��F� 9�j�]�o�����ğ�� �۟����o��@���1��PN�m�r� �mP��������P̯ ���`�*�/�� f`J�i�n�惹`����<���V 1���ށ��@]s8��T?HR_INRA �q�]مd�MASS6)� Z=�MN(�[��MON_QUEUE ������!UބN*�Un�Nk��ȫ�END��Ώ���EXE�����pBE����ϫ�OPTIO���׋��PROGR�AM %��%��習��TASK�_It �OCFG� ��π�ߵ�D�ATAx����G2�$�6�H�Z�l� ������������� �2���INFO
x�혝������ ����������	- ?Qcu��������N�Z��� �����pK_��ѳ��z�5G��2��D X,		�x�=���'�@���$a�����0_EDIT �������WERFL��Ó#�RGADJ �&�AЛ@R$?�]%�0�5&��?�����?���A<��z�%�o�/)(/�s#2�'"	Hʥ�l�!?8w�Aٴ�t$26�*A0/C2 **:L2�??Q3m=���2�5��+1�9��/�?y=�=�?�? �?�?�?KO�?O5O+O =O�OaOsO�O�O�O#_ �O�O___�_9_K_ y_o_�_�_�_�_�_�_ �_goo#oQoGoYo�o }o�o�o�o�o?�o�o )1�Ug�� ������	��� -�?�m�c�u���� ُϏ�[���E�;� M�ǟq���������3� ݟ���%���I�[� ��������ǯ������	�ߖ�𰄿�� ��39߿53��ϧ�0��B�o'PREF ��*00
5%I�ORITY:���>9!MPDSP8�'*��"��UT��34&OoDUCT����E��&OG_T�G$ �����TOE�NT 1�� �(!AF_IN�E��Y�J�!t�cpdߌ�!u�d{ߴ�!ic�m���.��XYx#�v��1)� Y1�*�0��S�6� B��f�������� ����!�3��W�>�{���*��x#�)�"�/X������Y7/c<H��44��(�.A�"?,  �u�(�}���+%�^Ŀ�f�x�,9!PORT�_NUM��0��9!_CART�REP% �aSK�STA�� 4L�GSV������#0Unothing����L��]TEMP �����T��_a_?seiban�,/ �</b/M/�/q/�/�/ �/�/�/�/�/(??L? 7?p?[?�??�?�?�? �?�?O�?6O!OZOEO WO�O{O�O�O�O�O�O �O_2__V_A_z_e_ �_�_�_�_�_�_�_o>�VERSI�����M` dis�abled'oSA�VE ���	�2670H782J�o�o!$�o�o���o 	x��V��	.�eKt���J�c|�o���mb]_� 1����`*�p�!�4�F��W��URGE_ENB�Ъ�(���WFr�DO���+�WRГ����WRUP_DE?LAY �,���R_HOT %�{���#���R_NORMAL����<W�&�SEMI6�\�|��U�QSKIP�	��#�xo��	o� �(���Y�G�}��� ��g�ů��կ���� �C�1�g�y���Q��� �������	�Ͽ-�� =�c�uχ�Mϫϙ��� ���Ϲ��)��M�_��q����$RBTI�F��0RCVTMkOUE�����DCR�Ǿ� ����C04^�@����3���띭3���*{vJ��-�7����I�4�<�	<�S�;�9<���<#*o<��M�Q 7���y��������/��A�S�e�w������R�DIO_TYPE�  ����EFPOS1 1�ui� xA
-���G 2k�o�*�N� ���1�Ug N���n� �/�/Q/�u// �/4/�/�/j/|/�/? ?;?�/_?�/�??�? �?T?�?x?O�?%O7O��?�?OOjO�O��O_S2 1�ԋ�ZO�O_�O6_�O��3 1��O�O�O,_�_��_�_L_S4 1� c_u_�_�_?o*oco�_S5 1��_
oo�Vo�o�o�ovoS6 1͍o�o�o�oiT|�S7 1�"�4F���"��S8 1Ϸ����~���5�SMAS/K 1���  ��� �ՇXNO���x:�D���MOTE���=�Z�_CFG ��a���A���PL_RANG]��ߛ�OWER �%��ΐ��SM_DRYPRG %%��%^��ԕTART� �ƞ�UME_PRO���p�=��_EXEC_EN�B  ���GS�PDI������Ѣ�T3DB����RMϯ���IA_OPTIO�N������U�MTE_݀T��_���*�fz��9���C�ˀ�����������OBOT_ISOKLC"�����ֵNAME %��_���OB_OR�D_NUM ?�Ƙ��H7�82  ˄h�@�h�$�hʬ�h�>�P?C_TIME�םٽx��S232z�1�����LTE�ACH PENDcAN��v�A�~��]�H@Maint�enance C�ons˂��ˆ"��DDNo Use~�E��i�{ߍߟ�8�ߵ���NPO#����A�!���CH_�LL��U���	�3���!UD1:�Y� �R܀VAIL�I����U�SRW  %������R_INTVAL����������V_DATA_GRP 2�%���X�D��P��W���{� f�%������������� ��$&8n\ ������� �4"XF|j� ������// B/0/R/x/f/�/�/�/ �/�/�/�/�/?>?,? b?P?�?t?�?�?�?�? �?O�?(OOLO:O\O ^OpO�O�O�O�O�O�O�_ _"_H_6_l_U���$SAF_DO_PULS��V���X���Q�PCAN������SC���(�����ˀq�����x�C�C��˂  p�o0oBoTofoxoo��o�o�o�o�o�o������be�!r �d�t:ql�(s�� @��fx��~Ny�� D�t�_ @�T�������T D�� *�S�e�w��������� я�����+�=�O��a�s�����`u2���ǟі��C�^��;�o2����p����
�t���Di���aC��  � ���Cђa x��Qa�s��������� ͯ߯���'�9�K� ]�o���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ�����������1�2��aZ�l� ~ߐߢߴ�������9� u�(�:�L�^�p��@�������2�0� D��N�	��-�?�Q� c�u������������� ��);M_q ������� %7I[m� ����D��/!/ 3/E/W/i/{/�/�/
� �/�/�/�/??/?A? S?������r�?�?�? �?�?�?�?O#O5OGO YOgIzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_�oo*o<oNo`o5�� ��9�ko�o�o�o�o�o &8J\n� ����pj�o�\�2���S�����	12345�678+�h!B�!ܺ�4���`��|�������ď ֏������o5�G� Y�k�}�������şן �����1�C�U�f� $���������ѯ��� ��+�=�O�a�s��� ����h�z�߿��� '�9�K�]�oρϓϥ� ���������Ͼ�#�5� G�Y�k�}ߏߡ߳��� ��������1�C�U� �y���������� ��	��-�?�Q�c�u� ������j������� );M_q�� �������% 7I[m��� ����/!/3/E/ W/{/�/�/�/�/�/ �/�/??/?A?S?e? w?�?�?�?�sm��?��?q/OO*OF��Cz  Bpqj �  ��h2�b�m�} ph
�G_�  	��r2�?`�O�O�O�Ook>�_D	lo�<��OB_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o'_�o�o�o�o (:L^p��� ���� ��$�>I�SB�1�AiB<S���$SCR_GR�P 1��8�� � � }�SA dE�	 ����������1B����SG��ۏɏ�:Mi�s@��D^@D/^�E��� \AR�C Mate 1�00iD/145�0ҁAM�ҁ�MD45 678�SC
12345��9��ӅE����KyBד_��SF�߃�@ S��Ó��Ӂ�	yJ�6�H�Z�l�~�SD���H������ ���Əǯ���Ά�oSAگC�֯g�N���v�B�M@Ʋ���ɴr��A^@ؿ  @S@�𵬁@��� ?PŬ�HM@)�ۺ��F@ F�`S� [�~��jϣώϳ��� ������!ߤ�� �L�07�I�[�m�B�{�� �߬�����	����?� *�c�N��r��_�� )������dG�@���0�SB�@P6���6�J����p�M@�������߃�?���SDA�������$�� QƒSA 3E��!ht�U (� ������� �$SF_�E�L_DEFAUL�T  ����S@@HO�TSTRL��`M�IPOWERFL�  BEX?�W�FDOM �R�VENT 1������w L!�DUM_EIP�.���j!AF�_INEL/SD!'FT�@./d/9!���/ �S/�/�!RPC_MAIN�/�(��/�/�#'VIS�/�)��/H?o!TP;0PU??��d7?�?!
PM�ON_PROXY�?�e�?�?[2�?��f�?,O!RDMO_SRV-O�gO�xO!R���O�h,gO�O!
� M�?��i�O_!RLSgYNC_��8�O>\_!ROS��\��4K_�_!
CE>]0MTCOM�_��k�_�_!	�RCO�NS�_�l�_@o!}�RWASRCGO��m/o�o!�RUSB�o�n{o�ow/ �o;C�o�o%Jn�5�Y�:RVI�CE_KL ?%�� (%SVCPRG1����u2�
��p3-�2��p4U�Z��p5}����p6�����p7͏ҏ�pH����9�"��t �OJ��q�r��q��� �qG��qo���q�� ��q��:��q�b��q ����q7����`�گ �������*��؟ R�� �z��(���� P�ʿ�x������ �ȯB�D����r�p ��p����<������� �	�B�-�f�Qߊߜ� ���߫��������,� �>�b�M��q��� ��������(��L� 7�p�[���������� ������6!Zl W�{�������2V�z_D�EV ���MC:��T4���pGRP 2������pbx 	� 
 ,�^����/�&/ //\/C/�/g/�/�/ �/�/�/�/?�/4?? X?j?��?E?�?�?�? �?�?OOOBO)OfO MO_O�O�O�O�O�O�O �O_q?_P__t_[_ �_�_�_�_�_�_o�_ (ooLo^oEo�oio�o �o�o�o3_ �o6 ZAS�w�� �����2�D�+� h�O������oy�� ��ߏ��@�R�9�v� ]�������П����۟ �*��N���C���;� ����̯ޯů��&� 8��\�C�����y��� ��ڿ��ӿ�g�4�F� -�j�Qώ�uχ��ϫ� �������B�)�f� x�_ߜ߃�����)��� ���,��P�7�t�� m����������� (��L�^�E�����w� ��o����� ��6 ZlS�w�� ����D��d Ԗ�	2{f������O%�x�/�����4! �4%D/R'</r/`/�/ �/�/�)/�/0)�/? ?>?,?N?P?b?�?�/ �?�/�?�?�?OO:O (OJO�?�?�O�?pO�O �O�O�O_ _6_xO]_ �O&_�_"_�_�_�_�_ �_oP_5ot_�_hoVo �ozo�o�o�o�o(o Lo�o@.dR�v �� �$��� <�*�`�N�������� t���p�ޏ��8�&� \�����L�����Ɵ ȟڟ���4�v�[��� $���|�����¯į֯ �N�3�r���f�T��� x��������:��J� �>�,�b�Pφ�tϪ� ���Ϛ�ߖ��:� (�^�L߂��ϩ���r� ���� ����6�$�Z� �߁���J������� �����2�t�Y���"� ��z�����������:� 1��
��R�v ����6�* :<N�r�� ��/�&//6/ 8/J/�/��/�p/�/ �/�/�/"??2?�/�/ ?�/X?�?�?�?�?�? �?O`?EO�?OxO
O �O�O�O�O�O�O8O_ \O�OP_>_t_b_�_�_ �_�__�_4_�_(oo Lo:opo^o�o�o�_�o o�o �o$H6 l�o��\~X� �� ��D��k�� 4������������ �^�C����v�d��� ����������6��Z� �N�<�r�`������� ��"��2�̯&��J� 8�n�\���ԯ������ �~���"��F�4�j� ����пZ��ϲ����� ����B߄�iߨ�2� �ߊ��߮�������� \�A��
�t�b��� �����"������� ��:�p�^��������� ����� "$6 lZ�������� �� 2h� ��X����
/ �/p�g/�@/�/ �/�/�/�/�/?H/-? l/�/`?�/p?�?�?�? �?�? ?OD?�?8O&O \OJOlO�O�O�O�?�O O�O_�O4_"_X_F_ h_�_�O�_�O~_�_�_ o�_0ooTo�_{o�o Dofo@o�o�o�o�o ,noS�o�t� �����F+�j �^�L���p������� ܏��B�̏6�$�Z� H�~�l����
�۟� �����2� �V�D�z� ������j�ԯf��
� ��.��R���y���B� ����п������*� l�Qϐ�τ�rϨϖ� �Ϻ����D�)�h��� \�J߀�nߤߒ���
� �����ߴ�"�X�F� |�j���������� ��
���T�B�x��� ����h��������� P��w��@� �����X~ O�(�p��� ��0/T�H/� X/~/l/�/�/�//�/ ,/�/ ??D?2?T?z? h?�?�/�??�?�?�? O
O@O.OPOvO�?�O �?fO�O�O�O�O__ <_~Oc_u_,_N_(_�_ �_�_�_�_oV_;oz_ ono\o~o�o�o�o�o �o.oRo�oF4j Xz|���* ���B�0�f�T�v� ��Ï������� �>�,�b�����ȏR� ��N�̟�����:� |�a���*��������� ȯ�ܯ�T�9�x�� l�Z���~�����Ŀ� ,��P�ڿD�2�h�V� ��zϰ�����Ϡ��� ��
�@�.�d�R߈��� ����x���������� <�*�`�߇���P�� �����������8�z� _���(����������� ����@�f�7v�j X�|���� <�0�@fT� x����/� ,//</b/P/�/��/ �v/�/�/?�/(?? 8?^?�/�?�/N?�?�? �?�? O�?$Of?KO]O O6OO~O�O�O�O�O �O>O#_bO�OV_D_f_ h_z_�_�_�__�_:_ �_.ooRo@obodovo �o�_�oo�o�o* N<^�o�o��o �����&��J� �q��:���6���ڏ ȏ���"�d�I���� |�j�������֟ğ�� <�!�`��T�B�x�f� ������ү���8�¯ ,��P�>�t�b���گ ��ѿ�������(�� L�:�pϲ���ֿ`��� ��������$��Hߊ� o߮�8ߢߐ��ߴ��� ���� �b�G���z� h��������(�N� �^���R�@�v�d��� ���� ���$����� (N<r`���� �����$J 8n���^�� ��/� /F/�m/ �6/�/�/�/�/�/�/ ?N/3?E?�/?�/f? �?�?�?�?�?&?OJ?�L1�$SERV_MAIL  T5�J@�0HOUTP�UT?H�0HRV 2��6  M@ (�1O�O�4DTOP10 2}�I d P? �O�O__/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o�������5�EYPE�`LNEFZN_CF�G ��5�MCL4oB�GRP �2�%�� ,B�   Ae�L1D;� Bf��  �B4L3RB2�1�FHELL�!��5��@�O<�Ώ>K%RSRݏޏ ��)��M�8�q�\��� ����˟���ڟ����7�I�[��  ��+�[�����i��� L0��ŢơL8q��2L0d�������H�K 1瞋  ˯@�J�D�n������� ��߿ڿ���'�"�4��F�o�j�|ώϊ�OM�M 螏�Ϗ�FTOV_ENB?D��A��OW_RE�G_UI��2BIM�IOFWDL���x��h�3�WAIT��A��oE^�Z@��D�X�TIM���ƒ�VA>@i�3�_U�NIT�����LC��TRY���4@MON_ALI_AS ?e���@heOM�_�q��J ;���������� � 2�D�V��z������� ��m�����
.�� Rdv�3��� ���*<N` �����w� //&/8/�\/n/�/ �/=/�/�/�/�/�/�/ "?4?F?X?j??�?�? �?�?�?�?�?OO0O �?AOfOxO�O�OGO�O �O�O�O_�O,_>_P_ b_t__�_�_�_�_�_ �_oo(o:o�_^opo �o�o�oQo�o�o�o  �o6HZl~) ������� � 2�D��h�z������� [�ԏ���
��Ǐ@� R�d�v���3�����П ⟍���*�<�N��� r���������e�ޯ� ��&�ѯJ�\�n��� +�����ȿڿ쿗�� "�4�F�X��|ώϠ� ����o�������0� ��T�f�xߊ�5߮��� �����ߡ��,�>�P��b���$SMON�_DEFPROG &������ &*SYSTEM*i�~���<{��RECALL ?�}�� ( �}�����
��.�@�R�  ��w�����������d� ��+=O��s �����`� '9K�o�� ���\��/#/ 5/G/�k/}/�/�/�/ �/X/�/�/??1?C? �/g?y?�?�?�?�?�? f?�?	OO-O?OQO�? uO�O�O�O�O�ObO�O __)_;_M_�Oq_�_ �_�_�_�_^_�_oo %o7oIo�_moo�o�o �o�oZo�o�o!3 E�oi{���� V����/�A�S� �w���������яd� ����+�=�O��s� ��������͟`��� �'�9�K�ޟo����� ����ɯ\�����#� 5�G�گk�}������� ſX������1�C� ֿg�yϋϝϯ����� f���	��-�?�Q����+copy mc�:diocfgs�v.io md:�=>192.16�8.56.1:17836Tߤ߶������5h�frs:o�rderfil.�dat virt:\temp\ߠ��,�>�P���-��*.d�����������xyzrat?e 124 t�� ��)�;�M������������������8�����mpback� ���.@R }/h�dbp�*��������3x��:\q� �� �-?Q��4�a�� ��������� ,/>/P/c��/�/��/�/���$SNP�X_ASG 2������!��  0��%y��/?  ?��&�PARAM ���%�! �	*	;P������o4��� OFT_K�B_CFG  ����%�#OPIN_�SIM  �+�j2�?�?�?�3� R�VNORDY_DOO  t5�5B�QSTP_DSB�>j2HO�+SR ���) � &�n:�O���&TOP_ON_ERRO~�FPTN �%��@�C�BRING_PRM�O�#BVCNT_GP� 2��%l1 0x 	DO?_��-_f_Q_�_�'VDPRP 1�C9m0{Q�1m_ �_�_�_�_o4o1oCo Uogoyo�o�o�o�o�o �o�o	-?Qc u������� ��)�;�M�_����� ������ˏݏ��� %�L�I�[�m������ ��ǟٟ���!�3� E�W�i�{�������د կ�����/�A�S� e�w���������ѿ� ����+�=�d�a�s� �ϗϩϻ�������� *�'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ����������1�C� U�|�y����������� ����	B?Qc�u���RPRG_�COUNT�6��B�	ENB�O�M���4�_UPD �1�nKT  
 �Y"ASe��� �����//+/ =/f/a/s/�/�/�/�/ �/�/�/??>?9?K? ]?�?�?�?�?�?�?�? �?OO#O5O^OYOkO }O�O�O�O�O�O�O�O _6_1_C_U_~_y_�_ �_�_�_�_�_o	oo -oVoQocouo�o�o�o �o�o�o�o.); Mvq����� ����%�N�I�[� m���������ޏُ���_INFO 1Y�/ �� � R�=�v�a��������YSDEBUG� �0���d��SP�_PASS�B�?�LOG �v/9  ��9���  ���UD1:\�<ϟ �_MPC$�/H����/[�Я /~��SAV �'�`���G�_���f��SVԛTEM_T�IME 1�'��: 0үf�ўT�SKMEM  t/�G�  ���%s���Ͽ��� @���� �������)U��A������TJ�\�n�(���� �Ϧϸ���^��'� W����p�+� =�O�a�s߅ߗߩ߻� ��������u�9� K�]�o������� �������#�5�G�Y��k�}���T1SV�GUNS*�'����ASK_OPTION� /:���_DI�����BC2_GRP� 2�/�Q���@��  C�:��BCCFG ��� ����` ��������! E0iT�x� ����/�/// ?/e/P/�/t/�/�/�/�/�/?���,!?�/ T?f?�/C?�?�?�?�? �?׮O���0O2O O VODOzOhO�O�O�O�O �O�O�O_
_@_._d_ R_t_�_�_�_�_�_�_ o�_oo*o`oFh10 to�o�o�o�oFo�o�o �o"FXj8� |������� 0��T�B�x�f����� ��ҏ�������>� ,�N�P�b�������ro ԟ���(���L�:� \���p�����ʯ��� ܯ� �6�$�F�H�Z� ��~�����ؿƿ��� �2� �V�D�z�hϞ� �Ϯϰ��������ҟ 4�F�d�v߈�߬ߚ� ��������*���N� <�r�`������ ������8�&�\�J� l��������������� ��"XF|2� �����f� B0fx�X� �����/// P/>/t/b/�/�/�/�/ �/�/�/??:?(?^? L?n?p?�?�?�?�?� �?O$O6OHO�?lOZO |O�O�O�O�O�O�O_ �O2_ _V_D_f_h_z_ �_�_�_�_�_�_o
o ,oRo@ovodo�o�o�o �o�o�o�o<�? Tf���&�� ���&�8�J��n� \���������Əȏڏ ���4�"�X�F�|�j� ������֟ğ���� �.�0�B�x�f���R ��Ư������,���<�b�P���p���A���*SYSTEM�*��V9.005�5 ��1/31/�2017 A �v  ��K�T�BCSG_GRP�_T   \ �$ENABLE��$APPRC�_SCL   
$OPEN��CLOSE�S_�MINF2'�AC�C��PARAM�� ���MC_MAX_TRQ�{$d�_MGNk��C�AVw�STA�Lw�BRKw�NO�LDw�SHORT?MO_LIM�ʧ�rh�J����PL1��T6���3��4��5���6��7��8k������� )$D�E�E��T��b�PATH^�w�m�~w�_RATIOk��s�T� 2 	/$CNT�A������m�INX�_UC�A���CAT_�UM��YC_ID� 	����_E�����6������PA�YLOA��J2L�_UPR_ANG6�LWA�?�3�O�x��R_F2LSHRTv�LOD���}��������ACRL_S��ؽ���+�k�HVA��$Hx���FLkEX�B�J2�w P�B_F��{$��_FTM���&��$RES�ERV�>�;��� ���� ;:$��LEN.�z�;�DE|���;�Yғ�����SLOW_A{XI��$F1��I��2��1�������MOVE_TIM���_INERTI���
�	$DTORQUEX�3��#}I��ACEMN��P%E�%Ep	V���d�A�R�TCV ��Rt����
��ET@�RJ���	M��,��J_MOD������ dRy�2��PpE���\�X��AW�gQ�JK@��K��V�K�VK�JJ0l���JJ�JJ��AA��AA�AA�%�AA �t�N1��N �d�#��E_�NU��A�JCF�G� � $�GROUPc�SK���B_CON�C���B_REQUI�RE���BU��U/PDATT�EL}  �%� �$TJ��� J�E��CTR��
T�N F�&�'HAN�D_VB��O�P� $oF2�x�3�m�COMP_�SW��@�R��O $$Ma�e�R�À�8���<� �5�¼6AI_.�h�D�<q�A��A��A��A���0��UD��D��D��P��3GR�ǂAST�ǂA4�ɂAN��DY��� x��4�5A���s��s� ��2�B��R����P����� �)�2�8;҆#� �0i�\� 7�U6��QA'SYM��
�TС���мݎ���_SH �"�������TU8����%�7�J>���P�pc�fio�_VI83��h6þ`V_UNI���d�{�JU�bU �b���d���d v��@��������su���x ���HR_T���	N2�q���DI�����O�te�p�#S
  �2I�QAz� ���q �S�s � B�� �p  � -f1MEe���4pr�QT�pPT&`r a�>���~$�5`C��^�R�T4`! $DUMMY1��$PS_ RF���$����FLA� YP_��F�$GLB_T�0 �u΅>���B�; 1�q� X��'�ST�f� SBRv�M�21_VT$S/V_ERa�O(`��,�CL��Ap Ol�r�pGL�`EW걿 4 $H�+$Y�2Z�2Ww���x�b3A���@�Y�U.]� oN��)`�$GI0}$>]� W����� Lh���'b}�$F'bE��NEA�R_ N��F�\ T�ANC��@�JOG���� �q$J�OINT�& ��MwSET�  ��E�� S�✔�!���  U�e?�� LOCK�_FO��m1�pBG�LV3GL��TE�ST_XM�j�EMP=�Ϣ悖��$UC�\���2� ������i0������CE| Ó� �$KAR�M�sT�PDRA`�3�*�VcEC~�D�.�IU����!CHE��TOOiL��i�V��REK�'IS3;���6��ЧACHP���v�O���F���29���I���  @$RAIL_BOXE��� ROBOƤ?���HOWWAR���屖���ROLM ���q!��¡!Ӱ���J�O_F� ! �����K�6���RN�Oo�W���?��C�<2Y�OUR������Q�"�!��/$PIPǦN]��Ӳ�� ��V�@�CORDED����u��q�� O�p  D ̀OBA�#��������̀��'`�!S;YS��ADR�!�p�>�TCH�0 � ,oEN�r#�A���_��d�z!�%P�VWVA� Ǥ 9�]��uPR�EV_RTA$�EDIT��VSHWR�!�&��]q�%�`D(�.Q��6Q?$HEAD8amp4��Ha��KEq�|��CPSPD�JM�P�L�u �TR�a �t���\�IjРS�"C20NEr�<�!�'TICK���Q�M�! g�:�HN�� @�W�~%��_GP��ʶ$�S3TY^ү�LO�ڠ��:��� t 5
��Gj�%$�Ѳ�u=��S�!$�a Jp-����p��P�P��SQU-������aT�ERCB����TS�$ ����' ]�'-`�>pOC�6�FbPIZ���������PR������S��P9U�a��_DO�c��XSN�K�vAXI4��/���UR� p@�"찕�"�]1� _`�4�ET5P��ЦU%��F�W��A�A�Q��ĳ��!5�� {SRE4lu� �9��:��6�	�2� �7��9��9�G� G�'F"TIF �R&��4CE op2oDoVd�!SSCЀ�  h� DS���4���SP�p"%A	T@�2���c⅂�ADDRESs�B���SHIF�#�_W2CH� �It!�TU�I�1 �W�CUSTOTVs1V��I�r U�P��6!��P
Ϫ
F�qV������! \���������,��J�2C�SC��Y�*��2�1�TXSCREE���"�p�TINA�O���T4����j�Q9_6"vP# TI�/� ��4�.���63��4��RRO�@�3а
��1�&�UE?�$# ��PMѧ�SP�4��RSM����UNEaX_�vA�pS_���+F�SA.IIG�S6Cx��B�4 2#O0UErT%�r?�nF��WGMT3pL�a��O@���BBL_r��Wo���& ���j�BO���BLEf"��C밚"�DRIGH��CBRDA�\!CKsGRo�UTEX$ |UQWIDTH������Ʊ��Jq�0I�>�EY6 ��' d�h��Ѐ���Ӱ��B�ACK�ᡂ�UE��!�FO���WLAB��?(!�I����$UR��PU�_P'�}H�1 ( 8wqB�_��t"�R(�Rq�@���������1�POm!J��)��L�PU�@r7cR���LUM7c�V ERV���SP��fT*�j GE��R�a `�)�LP$�e_E\���)�g���h!�h���i5�k6
�k7�k8�bZ�6���P�4������SJ�)^QUSR]�'+ <��'�U���#涒FO� ��PRI�rm��%q�pTRI}Pϱm�UN�p
�t,����p������� ��3 -� q-�RSp��G  �aT/��u!�rOSF���vR9 �2�so���.�f�x�������U�a��/$�6�DC�b��N�sOFFŠ��0���L�O�� 1.h9�����/9�GU.сP��A�׃��sQS�UB��H��@SRT���1���;���O9R��'�RAU� (�9T=�Z��VC� Ҕ2� ɲ��$�A��y�8񹳬`C��^{�DRIV��@C_V�����Ѐ�D4t?MY_UBY3t������$��19�l0��8	����P_S��l���BM�A$b�7DEY_�EX�@�3\����_MU.�X�An� @USA8��p[�@k0w�xp� �2x�Gg�PACINr�!�RG�𦥽�����A���SCp�RE�Rj!o�b�q`���S�3 Y�/TARGÐP72�$h�a�R�S�4nP0`�TQ�	o���RE6z�SW��_A��d�Io���OIq\!An v��E$pU�෱d��)�HK��5�����W�s��0��EA��ɷWOR�Pv����MRCV�A6 U��`O��M�PC83�	����REF �G(����e�s`cM� Xp�^��^�-ˀ����_RCʻ���0S!pf�ϓ��U�)��D7 ���gPTU0 epԕw�OU�����枃� 2��2�`$U00��r�4�5#�^�K SUL6b�5c`CO�0 `6`�]��Ӥ0����@��a��@q��i�L����$���a��@q�|s�?�8| +5#�k� 5#CACH��LOR�&�<�a�A��KQC ��C_LIM-Ig#FRj�Tl�N��$HO�P�*�OCOMM��BO�@���ب �a��VPH��/ ��_����Z�����k���WA{�MP��FAIk�G���;�AD?�p�IMR1E�_���GP@V��� k�ASYNBU=Fk�VRTD����l��&SOLo D_|���WA�P�ETU�O�X�Q����ECCU�VEM٠%�k�VIRC?����|B��_DELA�����p�p�AG��R�c�XYZM@5Cc�W3�qsQ T���r\P�s��D9�"�QLAS�AP6�
�� Gl� :��rX�Sa�7�N�m��VLEXE�;Ȕ3W�ka5!��FL2PIW���FI����F����q9#
�<_p�
��8t@s\���@ORD|q����##�� =_0Z`T��r�B�OJP6b��VSFE �3> a a0s���c�UR��M�u?�rV�R �J� f��"�5q@�r��qLIN��6@�WN�XS屎 QA��2��K&SHd`�HOLk(�XV�R�tB��@T_O�VRk��ZABC�C��"q-1��Zހ�tD�rDBGKLV��Lϒ�R�1_ZMPCF�E�d0�t2ޑLN~ �6�
� Mc��F �Ђ`��ɰ4CMC�M��C��CART�_Y14�P_2` O$Jw3q4D��}2�2�7`�5`6�U9X|5UXEu��6|�5�4�5�1�1�9��1�6�AZ�%G �+�$ `AY�V D�p H�RRM�{q��HET���R�PU'�Q1P�I � �3�� �PEAKf���K_�SHI�B��'RVB F^`G½B� C�@ r2g1|�����A20���I S��DXTRA�CE�PVw��AS�PHER'aJ �,e�THjO|I��$�TBCSG� 2� ����Q�����0  
 ` �_�_�_ �_�_�_�_�_.ooRo�dkwR~S�\d� ��a?�Q	 �HCBdo�iC  B �R�o�h�o�k#B��op��o�j9df  AXp? �w{qW�{������@�@0:nT� g�z�E�W���������
���3�	�V3.00�R	�md45�	*�U�M����1�� q��m���  ��X֟�wQJ2{c�]p6����  �U��Q ����rE�şp��p�����	_�ȯ���ׯ ���4��D�j�U��� y�����ֿ������� 0��T�?�x�cϜχ� ���Ͻ�������>�P�X�7�j�|�&ߜ� �߬�����	���-�� Q�c�u��B���� �������U%�7��Q ��=�c�Q���u����� ����������)M ;q_����� ��7%GI [������ ���//�M/;/]/ �/q/�/�/�/�/�/? ?%?�/I?7?m?[?}? �?�?�?�?�?�?�?!O OEO3OiOWOyO�O�O �O�O�O�O_�O__ /_e_S_�_w_�_�_�_ �_�_o�_+ooOo=o so�o//�o�o5/ko�o �o9'Io] ���u���� �5�G�Y�k�%���}� �������׏���1� �U�C�e���y����� ӟ������	��Q� ?�u�c���������ͯ ����o�oA�S��� +�q�������ݿ˿� �%�7�I�[���m� �ϑϣ���������� 3�!�W�E�{�iߋߍ� ������������A� /�Q�w�e����� ���������=�+�a� O���s�����e����� ����'K9[] o������� #G5k}�� [�����// C/1/g/U/w/y/�/�/ �/�/�/	?�/-??=? c?Q?�?u?�?�?�?�? �?�?�?)OOMO_O�� wO�O3OaO�O�O�O�O __7_%_G_m__�_ O_�_�_�_�_�_o!o 3oEo�_ioWo�o{o�o �o�o�o�o�o/ SAcew��� �����)�O�=� s�a���������ˏ� �O	��-�׏]�K��� o�������۟ɟ��� #�5��Y�G�}�k��� ��ůׯ������1� �U�C�y�g������� ӿ������	�?�-� O�Q�cϙχϽϫ��� ������;�)�_�M� �ߕ�?��߿�i���� ��%��I�7�m�[�}� ������������!�8�E�/�  e�i�� i�}�i��$�TBJOP_GR�P 21���  ?��i�	�������9� � ����� ���������i� @�e��	 �CB  ��C����5�GU	i�C 2BH  A�/��D�,��bAB* q�$�7C�� ���c��d��i�A �EG+��a	�0��D/�D<Ky/@�//#/�/�/�� 	??�/�/T?f?%?o? a	�?�?�?�?�?�?�? O)OO!OOO�O[OO��O�O�O�O�O_g��i�1Q�E	V3�.00��md45��*[P��d�i_�tW G/� �G7� G?h �GG8 GO �Gd� Gz  �G�� G�| �G�: G�� �G�� G�t �G�2 G�� �Gݮ G�l �G�* G�� �HS�RF� �F@ F+� �FK  Fj` �F� F�Q � GX �R�Q^�� Gv G��ĨS�4 G��� G�� G�\� G� =L�_�=#�
]Ae��Js�Yokbi��oo�o��ESTPA�R�P]����HR��`ABLE 1	*��C`i��h�g ��di�g�hn i��h�p�g	�h
�h��h�ei��h�h8�hDa�cRDI�o���o!3EWu�tO��{����+��bS��� �z��� �"�4�F�X�j�|��� ����ğ֟����� 0�B���Āȏ���g�� l�~�����N`r���x�bi�NUM [ 1���	 �q� C`D`�b_CFG 
R����@��IMEBF_�TT�a�����`��V�ERBc������R� 1�k 8$f_i�d�� P���  ���%�7�I� [�m�ϑϣϵ����� �����!�3�|�W�i߀�ߍߟߵ�������A0�����MD3�E���� k�}��V_qI����INT������T1�#�5� Bp��O�a���_TC�������$�P����9�R�Q��Դ_L���@�˵�`MI_CH�AN�� ˵ nD_BGLVL��˵��aq ETHERA�D ?�e� ��`�����hq oROUT��!P��!#ASNM�ASK�˳�255.GS}���GS�`OOLOFS�_DI�P�%�	O�RQCTRL !޻7��o-T/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c?�s</�?�?�?�cPE?_DETAI���PGL_CONF�IG R�b����/cell/�$CID$/grp1�?4OFOXOjO|O2��
�O�O�O�O�O _�O%_7_I_[_m__ _�_�_�_�_�_�_�_ �_3oEoWoio{o�oo �o�o�o�o�o�o/ ASew�*�@�������}� O�a�s���������?я������*�<� N�`����������̟ ޟm���&�8�J�\� n���������ȯگ� {��"�4�F�X�j��� ������Ŀֿ����� �0�B�T�f�x�Ϝ� ���������υ��,� >�P�b�t߆�ߪ߼� ��������(�:�L� ^�p������������ ��@�U�ser View� "I}}1234?567890C�U� g�y�������. C����)�26����+=Oa����0�3 �������	h*��4�cu�� �����5R/ )/;/M/_/q/��/��6/�/�/�/??%?�/F?��7�/?�?�?@�?�?�?8?�?��8n? 3OEOWOiO{O�O�?�O��B lCamera4�*O�O@__)_;_M_+�E�O w_�_�^A��_�_�_�_�_o)  �F���O _oqo�o�o�o�o`_�o �oLo%7I[m�O��F�	�� ���%��oI�[�m� �������Ǐُ돒 �wQ��7�I�[�m�� ��8���ǟٟ$���� !�3�E�W����w+k� ����ɯۯ�����#� 5�G���k�}������� ſl��E�)Z��!�3� E�W�i���ϟϱ��� ��������/�ֿ�w m9��{ߍߟ߱����� |�����h�A�S�e� w���Bߤw!I2��� ����/�A���e�w� �����������������9��HZl~ ��I�������� 2DVhz	J	�E0 ����� /�3/E/W/�{/�/ �/�/�/�/|��@�K y/.?@?R?d?v?�?// �?�?�??�?OO*O <ONO�/�EBk�?�O�O �O�O�O�O�?_*_<_ �O`_r_�_�_�_�_aO ��{Q_oo*o<oNo `o_�o�o�o�_�o�o �o&�_�U��o r�����so� ��_8�J�\�n��� ��9�U��)�ޏ��� �&�8��\�n���ˏ ����ȟڟ������U 򻕟J�\�n������� K�ȯگ�7��"�4��F�X�j��   �������Ͽ�����)�;�M�_�   o�w��ϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������������c�  
�(�  荰( 	 ��;)_ M�q�������%��� ̹�j|���� ���/�Y6/H/ Z/�~/�/�/�/�/�/ /�/? ?g/D?V?h? z?�?�?�/�?�?�?-? 
OO.O@OROdO�?�? �O�O�OO�O�O__ *_<_�O`_r_�_�O�_ �_�_�_�_oI_&o8o Jo�_no�o�o�o�o�o o!o�o"ioFX j|���o��� /��0�B�T�f�� �������ҏ���� �,�s���b�t���͏ ����Ο����K�(� :�L���p��������� ʯ�� ��Y�6�H� Z�l�~���ׯ�ƿؿ �1�� �2�D�V�h� ���Ϟϰ��������� 
��.�u�R�d�v߽� �߬߾�������;�@ �#�5�G���� ��0fr�h:\tpgl\�robots\a�m100id\a�rc_mate_���_1450.xml�������������0�B�T�E��� Y�~������������� �� 2D[�Uz �������
 .@WQv�� �����//*/ </SM/r/�/�/�/�/ �/�/�/??&?8?O/ I?n?�?�?�?�?�?�? �?�?O"O4OK?EOjO |O�O�O�O�O�O�O�O __0_GOA_f_x_�_ �_�_�_�_�_�_oo�,o>n`��� |�k�<< i�?�>k�o>oyo�o �o�o�o�o�o�o5 -O}c���������1�?��$�TPGL_OUT?PUT I�I�_ a`i� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ���
���i�a`�6�2345?678901A�S� e�w�������?�>�ʯ ܯ� ��$���(�Z� l�~�����:�}��Կ ���
�ϴ�ƿR�d� vψϚϬ�DϺ����� ��*���8�`�r߄� �ߨ�@�R������� &�8���F�n���� ��N��������"�4� ����j�|��������� \�����0B�� Px����Xj �,>P�^ �����f�/@/(/:/L/�A�}\a��/�/�/�/�/�/�-@�co?#?ij ( 	 &�X?F?|?j? �?�?�?�?�?�?�?O OBO0OfOTO�OxO�O �O�O�O�O_�O,__�<_>_P_�_t_�_4�� _`xf�_�_�]�_o*o oNo`o.��_�o�o=o �o�o�o�o!o% W�oC��y�� 3����A�S�-� w����q���яk��� ���=�����s��� �����������a� '�9�ӟ%�o�I�[��� �������ٯ#�5� �Y�k�ɯS�����M� ׿�ÿ��}��U� g�ϋϝ�wω���1� C�	�ߵ�'�Q�+�=� �ߙ��ϝ���i߻�� ���;�M��5��� o��������_��� 7�I���m��Y����� �%�������3 i{����K�����/�R�$�TPOFF_LI�M �P��Q���JN_SV�N  �$`P_MON �USb��2�%�JSTRTCHK' �U`/h�VTCOMPAT�u�dVWVAR� �"(y K� :/Y��J_DEFPR�OG %�%�Q/�/f_DISP�LAYU�j"IN�ST_MSK  �, �*INU�SER��$LCK��,�+QUICKM�EN"?�$SCRE�A0�U "tpsc�$�!\0a9`�r0_v9ST�`R�ACE_CFG ��"$Y	�C$
?��8HNL� 2y*�P�1)+  O"O'O9OKO]OoO�O��O�J�5ITEM �2K �%$�12345678�90�O�E  =<��O_*_2S  !8_@[L �O�_C#�O �_
_�_�_@_�_d_v_ ?o�_Zo�_jo�ooo o*oDoNo�oroD V�oz�o�o|& ��
�n���� :��������"�ʏF� X�!�|�<���`�r�֏ ����L�՟0��T� � &�8���D���ҟ�^� ���گ�P��t��� ���4�ί������� (�:��^�ς�B�T� ��j�ܿ����6� ��ߎ�~ϐϢϼ��� @��ϖ߼���2���V� h�z��ߞ�J�p���� ��
��.�� �d�$� 6���B��������� �����N� r���M ��h��x��� 8J\��,Rd ������F //|$/��{/� �/��/�/0/�/T/f/�/?�4S�2�?4:ψ  �B4: 8�1�?�)
 �?�?��?�?c:UD1:�\�<��F1R_G�RP 1�K?� 	 @� :O LK6OlOZO�O~O�O�N��@�O�J�A�?_�O<7_"U?�  R_d[ N_�_r_�_�_�_�_�_ �_�_&ooJo8ono\o0�o�o�o�o	5�o��oD3SCB 2P; =_:L^�p�����:<U�TORIAL �P;�?�?7V_C�ONFIG  �P=�1�?�?t�$�OUTPUT !P9e�����ď֏ �����0�B�T�f� x�����b���ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϷ� ������ ��$�6�H� Z�l�~ߐߢ߳����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� �����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/N�`��� �/??&?8?J?\?n? �?�?�?�?�?��?�? O"O4OFOXOjO|O�O �O�O�O�?�O�O__ 0_B_T_f_x_�_�_�_ �_�_�O�_oo,o>o Poboto�o�o�o�o�o �_�o(:L^ p������o�  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�nπ�ϒϤ϶����Ͻ(���������� 6��/Z�l�~ߐߢߴ� ��������� �2�� V�h�z�������� ����
��.�@�Q�d� v��������������� *<M�`r� ������ &8I\n��� �����/"/4/ F/Wj/|/�/�/�/�/ �/�/�/??0?B?S/ f?x?�?�?�?�?�?�? �?OO,O>OO?bOtO �O�O�O�O�O�O�O_ _(_:_L_]Op_�_�_ �_�_�_�_�_ oo$o 6oHoY_lo~o�o�o�o �o�o�o�o 2D�S{�$TX_SCREEN 1"�����}�S�������Bք1�C�U�g� y�������ӏ��� 	����?���c�u��� ������4��X��� )�;�M�_�֟蟕��� ��˯ݯ�f����7� I�[�m�������,� ٿ����!�3Ϫ��� i�{ύϟϱ���:��� ^���/�A�S�e�������$UALRM_MSG ?sy��p ��Vj���� ����"��F�9�K�i�o���������S�EV  ������ECFG �$su}q  �Ve@�  AJ� �  B�Vd
  ��]csu}��������� ������1?&�GRP 2%0�; 0Vf	 g�����I_BBL_N�OTE &0�T��l]b�xp_a<�DEF�PRO��Z�� (%��_`�* N9r]�������/�FKE�YDATA 1'<sys p ?�Vf =x/�/� g/�/�/�%,(/�/Vd �/??C?*?g?y?`? �?�?�?�?�?�?�?O -OOQO8OuO�OnO�O �O�O�O�O_�O)_X.��9_`_r_�_�_�_ �_]bN_�_�_oo+o =o�_aoso�o�o�o�o Jo�o�o'9K �oo�����X ���#�5�G��k� }�������ŏ׏f��� ��1�C�U��y��� ������ӟb���	�� -�?�Q�c�򟇯���� ��ϯ�p���)�;� M�_��������˿ ݿ�~��%�7�I�[� m�D_�ϣϵ������� ��!�3�E�W�i�{� 
ߟ߱��������߈� �/�A�S�e�w��� ������������+� =�O�a�s�������� ��������'9K ]o��"��� ���5GYk }������ //�C/U/g/y/�/ �/,/�/�/�/�/	?? �/??Q?c?u?�?�?�?ڂ��;�������?�?�=�? O2OF,_cO_�OnO �O�O�O�O�O__�O ;_"___q_X_�_|_�_ �_�_�_�_o�_7oIo 0omoTo�o�o���o�o �o�o!0?EWi {���@��� ��/��S�e�w��� ����<�я����� +�=�̏a�s������� ��J�ߟ���'�9� ȟ]�o���������ɯ X�����#�5�G�֯ k�}�������ſT�� ����1�C�U��y� �ϝϯ�����b���	� �-�?�Q���u߇ߙ� �߽����߸o��)� ;�M�_�f߃���� ������~��%�7�I� [�m������������ ��z�!3EWi {
������ �/ASew ������/� +/=/O/a/s/�//�/ �/�/�/�/?�/'?9? K?]?o?�?�?"?�?�? �?�?�?O�?5OGOYO kO}O�OO�O�O�O�O��O__��![�>�����J_\_ n]F_�_�_|V,�o�_ �o�_�_o-ooQo8o uo�ono�o�o�o�o�o �o);"_F� j������� ��7�I�[�m�����O ��Ǐُ����!��� E�W�i�{�����.�ß ՟�������A�S� e�w�������<�ѯ� ����+���O�a�s� ������8�Ϳ߿�� �'�9�ȿ]�oρϓ� �Ϸ�F��������#� 5���Y�k�}ߏߡ߳� ��T�������1�C� ��g�y������P� ����	��-�?�Q�(� u��������������� );M_��� �����l %7I[��� ����z/!/3/ E/W/i/��/�/�/�/ �/�/v/??/?A?S? e?w??�?�?�?�?�? �?�?O+O=OOOaOsO O�O�O�O�O�O�O_ �O'_9_K_]_o_�__ �_�_�_�_�_�_�_#o�5oGoYoko}o�of���k�f�����o�o�m�o �f,�C�gN�� �������� ?�Q�8�u�\������� Ϗ���ڏ�)��M� 4�q���b�����˟ݟ ��o%�7�I�[�m� ��� ���ǯٯ��� ���3�E�W�i�{��� ���ÿտ����� ��A�S�e�wωϛ�*� ���������ߨ�=� O�a�s߅ߗߩ�8��� ������'��K�]� o����4������� ���#�5���Y�k�}� ������B������� 1��Ugy�� ������	- ?Fcu���� �^�//)/;/M/ �q/�/�/�/�/�/Z/ �/??%?7?I?[?�/ ?�?�?�?�?�?h?�? O!O3OEOWO�?{O�O �O�O�O�O�OvO__ /_A_S_e_�O�_�_�_ �_�_�_r_oo+o=o Ooaosoo�o�o�o�o �o�o�o'9K] o�o��������� ��� ���*�<�N�&�p���\�,n���f�׏ ������1��U�g� N���r��������̟ 	���?�&�c�J��� ������������ )�;�M�_�q������ ��˿ݿ�ϐ�%�7� I�[�m��ϣϵ��� �����ό�!�3�E�W� i�{ߍ�߱������� ����/�A�S�e�w� ������������ ���=�O�a�s����� &����������� 9K]o���4 ����#�G Yk}��0�� ��//1/�U/g/ y/�/�/�/��/�/�/ 	??-???�/c?u?�? �?�?�?L?�?�?OO )O;O�?_OqO�O�O�O �O�OZO�O__%_7_ I_�Om__�_�_�_�_ V_�_�_o!o3oEoWo �_{o�o�o�o�o�odo �o/AS�ow ������r� �+�=�O�a������ ����͏ߏn���'��9�K�]�o�F q�}�F �����@���������̖,ޯ #�֯G�.�k�}�d��� ��ůׯ������1� �U�<�y���r����� ӿ����	��-��Q� c�B/�ϙϫϽ����� ����)�;�M�_�q�  ߕߧ߹�������~� �%�7�I�[�m��ߑ� ������������!� 3�E�W�i�{�
����� ����������/A Sew���� ���+=Oa s������ //�9/K/]/o/�/ �/"/�/�/�/�/�/? �/5?G?Y?k?}?�?�? x��?�?�?�?OO&? COUOgOyO�O�O�O>O �O�O�O	__-_�OQ_ c_u_�_�_�_:_�_�_ �_oo)o;o�__oqo �o�o�o�oHo�o�o %7�o[m� ���V���!� 3�E��i�{������� ÏR������/�A� S��w���������џ `�����+�=�O�ޟ s���������ͯ߯�0����0���
��.��P�b�<�,Nϓ�FϷ���ۿ �Կ���5�G�.�k� RϏϡψ��Ϭ����� ����C�*�g�y�`� �߄����߲?��	�� -�?�Q�`�u���� ������p���)�;� M�_������������ ��l�%7I[ m�������� z!3EWi� �������� ///A/S/e/w//�/ �/�/�/�/�/�/?+? =?O?a?s?�??�?�? �?�?�?O�?'O9OKO ]OoO�OO�O�O�O�O �O�O_��5_G_Y_k_ }_�_�O�_�_�_�_�_ oo�_CoUogoyo�o �o,o�o�o�o�o	 �o?Qcu��� :�����)�� M�_�q�������6�ˏ ݏ���%�7�Ə[� m��������D�ٟ� ���!�3�W�i�{� ������ïR����� �/�A�Яe�w����� ����N������+�h=�O�&PQ��&P���zόϞ�v����Ϭ�,��߶� '��K�]�D߁�hߥ� �ߞ����������5� �Y�k�R��v��� ���������1�C�"_ g�y���������п�� ��	-?Q��u �����^� );M�q�� ����l//%/ 7/I/[/�/�/�/�/ �/�/h/�/?!?3?E? W?i?�/�?�?�?�?�? �?v?OO/OAOSOeO �?�O�O�O�O�O�O�O �O_+_=_O_a_s__ �_�_�_�_�_�_�_o 'o9oKo]ooo�oX��o �o�o�o�o�oo#5 GYk}��� �����1�C�U� g�y��������ӏ� ��	����?�Q�c�u� ����(���ϟ��� ���;�M�_�q����� ��6�˯ݯ���%� ��I�[�m������2� ǿٿ����!�3�¿ W�i�{ύϟϱ�@��� ������/߾�S�e�@w߉ߛ߭߿ߖ`�����`�����������0�B��, .�s�&���~����� �����'��K�2�o� ��h������������� ��#
GY@}d ���o��� 1@�Ugy��� �P��	//-/?/ �c/u/�/�/�/�/L/ �/�/??)?;?M?�/ q?�?�?�?�?�?Z?�? OO%O7OIO�?mOO �O�O�O�O�OhO�O_ !_3_E_W_�O{_�_�_ �_�_�_d_�_oo/o AoSoeo�_�o�o�o�o �o�oro+=O a�o������ ���'�9�K�]�o� v������ɏۏ��� ��#�5�G�Y�k�}�� ����şן������ 1�C�U�g�y������ ��ӯ���	���-�?� Q�c�u��������Ͽ ���Ϧ�;�M�_� qσϕ�$Ϲ������� �ߢ�7�I�[�m�� �ߣ�2���������� !��E�W�i�{��� .�����������/���$UI_INU�SER  ����P���  0�4�_M�ENHIST 1�(P�  �( ]����(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1o�������9 ����936��d v��)���� ��ASew ��*����/ /�=/O/a/s/�/�/ �/8/�/�/�/??'? �/K?]?o?�?�?�?�<�D1��D?�?�?OO )O;O>?_OqO�O�O�O �OHO�O�O__%_7_ �O�Om__�_�_�_�_ V_�_�_o!o3oEo�_ io{o�o�o�o�oRodo �o/AS�ow ������?�?� �+�=�O�a�d���� ����͏ߏn���'� 9�K�]�o��������� ɟ۟�|��#�5�G� Y�k���������ůׯ ������1�C�U�g� y��������ӿ��� ��-�?�Q�c�uχ� ���Ͻ�������ߔ� )�;�M�_�q߃ߕ�$� �����������7� I�[�m��� ���� �������!���E�W� i�{�����.������� ����Sew �������� +��as�� ��J��//'/ 9/�]/o/�/�/�/�/ F/X/�/�/?#?5?G? �/k?}?�?�?�?�?T?��?�?OO1OCO.���$UI_PAN�EDATA 1*����yA  	�}UO��O�O�O�O�O�O ) �O_8�OG_Y_k_}_ �_�__�_�_�_�_�_ ooCo*ogoyo`o�o��o�o�o�o�o1	� @r/_4FX j|��o�%_�� ���0�B��f�M� ��q��������ˏ� ��>�%�b�t�[���|��{C�۟��� �#�5���Y��}��� ����ůׯ>������ 1��U�g�N���r��� ��ӿ�̿	��-�?� ��ğuχϙϫϽ��� "���f��)�;�M�_� q߃��ϧߎ��߲��� ���%��I�[�B�� f������L�^�� !�3�E�W�i������ ����������� A(ew^��� ����+O 6s�������� �//h9/��]/o/ �/�/�/�//�/�/�/ ?�/5?G?.?k?R?�? v?�?�?�?�?�?OO ��UOgOyO�O�O�O O�OF/�O	__-_?_ Q_c_�O�_n_�_�_�_ �_�_o�_)o;o"o_o Fo�o�o|o�o,O>O�o %7I�om �O������d !��E�W�>�{�b��� ����Տ������/�0�S��o�o}�d��� ����ӟ���)��� �u�H�Z�l�~����� 	�Ư���ѯ� �� D�+�h�z�a�����¿�Կ�����x�c�k�$�UI_POSTY�PE  �e� 	 ��[�*�QUICKM_EN  9�H��^�,�RESTOR�E 1+�e  ��B�r�����ϑrm � )�;�M�_�q�ߕߧ� �����߀���%�7� I���V�h�z��ߵ��� �������!�3�E�W� i�{������������ ������Sew ��>���� �+=Oas( ����//'/ 9/�]/o/�/�/�/H/ �/�/�/�/?�?0? B?�/}?�?�?�?�?h? �?�?OO1OCO�?gO�yO�O�O�Oi�SCR�Ey�?~��u1sc��u2��D3�D4�D5�D6��D7�D8�A�CTAT5�� ���e"ʏUSER�@�O�BTL�@�Cks�C�T4�TU5�T6�T7�T8�Q�*�NDO_CFG� ,9�t�s�*�P�D-QgY�?None *�^P�_INFO 1-j�e`��0%�O ,o�xo[o>oo�oto �o�o�o�o�o!�EW:{b��QOFFSET 09�a�PC��XO�� ��/�&�8�e�\�n� �r�����ȏ����� +�"�4�F����ϒ���ⵟ
��ڟ�xUFR�AME  PD��V�QRTOL_A�BRT���s�EN�B��GRP 1�1�Ɋ�Cz  A�u�s��Qs����������ͯ߯��x�U�?��Q.�MSK  �B�a.�N��%�	i�%b���k�VC�MR[�27�{�#�R@	�Pfr�1: SC130EF2 *ݿ�PDe�����T&��5R@��Q?��@�p:��ȇ� ɟ5�?�IH`�rϟ�ı�ϴ��8��A�RB����RB B����RA#ի�Dߋ� h�7ߌ�w߰ߛ��߿� ��
�a���@�+�=�v��)ߚ�ISIO�NTMOU�B���U���R8SﳸS� j� FR:\���\�PA\�� �߀ MC�LO�G�   UD�1�EX5�RA'� B@ �� x�I�r���I����PC� � n6  ���IFu�%���`��Z�  =���PD	 J�}*�TRAIN_����ǐ  dPQp	�栲9�}(c� �W����� ��.2@Rdhv���_\�RE���:b�ʲ��LEXEr��;�{�Q1-e��VMPHAS/P��U�SЖ�RTD�_FILTER �2<�{ Ԓ�� ,�{/�/�/�/�/�/�/ �/??��i/N?`?r? �?�?�?�?�?�?�?���SHIFT�1=�{
 <��q�JO DU)OOO�O_OqO�O�O �O�O�O�O_<__%_�r_I_[_�__	L�IVE/SNAP�esvsfliv\.�_��� �pyU�P�Rmenu�_��_�_Woio@b	E��>XIO�EMO��?��� ��$WAIT?DINEND��+���dO?�"��g���oS��iTIM@���<|G�o^}�o�{�az/azN�hREL�E%!@��d�����a_ACT�P�K�E�� @d�ko���E��RDIS�PA��`V�_AXSR�p2A�b�����Vp_I�R  +&��  	��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i�{�������ÿ�տ�������XV�R�aB��$Z�ABCp1C�� ,N f�2ϵ�Z[IP��D�e�������ύ�MPCF__G 1Eٍ0J��=��S�FىX�`#� �c�߆�<90 �߻�S�|��ߠ�?�}������ S��$�z�8���� ���������@��
�4�M���G��|JÛ�YLINDK!�Hً Є� ,(  *������`���������� �� );M��p���{ ��� U6 ��lS�w������Y�2Iه]� �)�#/3,���\/@G/�/��/�/���!�A�c�SPHER/E 2Ju��*? z�/<?#?`?��/�? �?$�?k?Q?O�?&O O?\OnO�?�?�OO �O�O�O�OEO"_4_F_6M�ZZ/� ǘf