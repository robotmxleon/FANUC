��   :�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����FSAC_LS�T_T   8� $CLNT_�NAME !�$IP_ADDR�ESSB $AC�CN _LVL � $APPP  _  �$8 AO ? ���z�����o VERS�IONw�  �׋IR�TUALw�'DCEF\ � � �� ����ENABLE� ������LIST 1 �  @!�$,��)���(y L^������ �-/ /Q/$/u/H/Z/ �/~/�/�/�/�/�/? �/:? ?q?D?V?h?�? �?�?�?�?O�?7O
O OmO@O�OdO�O�O�O �O�O_�O3___U_ <_z_`_�_�_�_�_�_ �_�W