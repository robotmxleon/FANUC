��   b�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����CELLSET�_T   �w$GI_STY�SEL_P }7T  7ISO:iRibDiTRA�R�>�I_INI; �����bU9AR�TaRSRPNS�1Q234�5678�Q
TROBQACKSNO� �)�7�E�S �a�o�zU2 3 4 5 6 7 8awn&GINm'D�&��) %��)4%��)P%�̖)l%SN�{(OU���!7� OPTNAA�73�73.:B<;�}a6.:C<;CK;C�aI_DECSN�A�3R�3�TRY�1��4��4�PTHCN�8D�D�INCYC@HG��KD�TASKOK �{D�{D�7:�E� U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V�8�Tb@SEGq�Tp��T�@REQ� d�drG�:Mf�GJO_HFAUL�Xpd�dvgALE�  �g�c�g�cvgE� �H<�dvgNDBR�H�dgRGAB�Xtb~���CLMLIy@�   $�TYPESIND�EXS�$$CL�ASS  �S��lq����apVERSIONix�  ���}qIRTUAL�i{q'61�r��ƒp��q�t+ UP�0 �xSt�yle Sele?ct 	  ���r��uReq. /E�cho���Ac�k���Ini�tiat�p�r�"
�^�m������e	��
��  ��������:q�����χ�q)��Op�tion bit# A<��p�B��}C4�Decis��codY��Try�out mj�6�Path segh�_ntin.8�Ig��ycX�:�Task� OK��?�Man�ual opt.%r�A���B����C� decsn� ��$�Robot� interlo�7�@�\� isolQ�4�C��iM�@���ment<�)��������Ě}�statu�s=�	MH Fa�ult:����Al�er�1�C��p@r 1�z j�;�y����I�; LE_CO�MNT ?�y�   Չ�ѿ� ����*�<�N�`�r� �ϖϨϺ�������� �&�9�J�\�n߀ߒ� �߶����������"�����U��9r��Ŵ �  ��ENAB  ��:�������������ꮵMEN�U\��y��NAME� ?%��(%$* R�זb��P���t��� ������������+ O:s^p��� ��� $6 HZ�~���� ���/ /Y/D/}/ h/�/�/�/�/�/�/�/ ?
?C?.?@?R?d?v? �?�?�?�?�?�?�?O M