��   �A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A   �����
�WVAMP_�T   �$X1  $kX2AY@</�FC5  �$2ENBA $�DT  / _�R2 d EN�ABLEDnSC�HD_NUMA � xCFG5�� $GROU�P�$z ACCE�L@�G$MA?X_FREQ�2 �L�DWEL�D�EBUG�PRE;WSOUT��PULSEAS�HIFt 7TYP�4$USE_A�EF} 4$GD=O�  f0� r?�NpW�EAVE_TSK� �V�_GP��SUPPORT�_CFnCNVT_DONE p �}k}GRP #2r�� _� ��$� TIME1�o$2'EXT�� (1#&(MODE�_SW�CO3 S�WIT �/ PH�AX6  4 �� ECC$�T�ERMNnPE�AKno!AL � \ � �!I֑$�!N_VSTAR�#!r"ؾ�"�%�CY{CL42 
���/ � Tv"b $�CUR_REL_�� �!3WPR5� � 
$CEN� _RI3RADkIU�XI�z ] ZIMUT�i!$ELEVAOTIONg5� N��CONTINUO�e2q �MEXAC�=PE�S�6 � H~ �UENCyYA�ITUD4��2RIGHC�2L}EBL_ANG1 �OTF_�� 	�  $3A�bET��n�3C!$OR�GjHFBKjH��P���C��DLDW�HR�E�_�3�B�C ��D�B�C�@�D�A�CCHG�G	Q�F	Q�F	Q�FINC�G=Q�F�=Q�F=Q�F�AVCPYC� _T�\#�Y~PL#�@SY��H)@��UPD"0n��$$CLASS ? ����Q��x8 �P�PVERS�1��W  ����QIRTUAqL�_�Q0 2�X�� � ?��@�  HaDae �TWoio{o�o�o`)d�N 2 3k �Hf��uHe@O�Hi�oNc)a� � eG� E`��`9t�12  ������=�����4s ����jpYq��w�r��1��xat� �ujp`��i.�5t�8q�q2�b�t���
F�9x������ ��̏ҏ���Sb)a� w 23k
TDa�SI�8� ������0h�?m�'����l�D�����Ca ��l����k��� �2��D�V�h�z��l�FIGURE 8��o�v�Hal�f��� �����M�(�H��󀈯������Ŀֿ�T�CIR1�� Pd�}�0�~�h�z�D�Z�l���0�v˜�~������ ��$ߪjN� Hp��4q�Ȓ���@��ʖD�M`g�� ��������	��-�?�pQ�c�u`��� �q� �5) �ᐟN`���ᬟ���� ˟���M�_�q������������kTriangle�� z�h߾�M��Ɵ�� �������/ L�& ��g�n���	/ /-/?/Q/c/u/�}D Vhz��/�/�� 9?K?]?o?�?�?�?�?�?����� O�h�� O2ODOVOhOzO�O�O �O�O�O�O�O
__.[ �?._O"O�_�_�_�_ �_�_�_oo&o8oJo�\ono�mSCHEXTENB  =���ctSTATE ;2�k |o�o��o �gWPR �7�6�L}D�-�_?OTF 	8��@)0�q�q���v)��uAȫs�u@�  <#�
�?��|��mu_GP 2w| ���d�v�� ��я㏡+