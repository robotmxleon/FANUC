��   K�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_���$$C�LASS  ������D��D�VERSION�  ���/IRTUA�L-9LOOR� G��DD<x$p?�������k,  1 <D
wX������ Z)/;/Z�/o/�/@�/a/�/�/�/_ �/��/	?';�$MNU�>A�  <���d?/\?~?�? �?�?�?�?�?O�?O 2O`O*cO�OwO�O�O �O�O�O_�O_E_�~;5NUM  ������PtUTOOLC?\ 
Y?[_�_ CO�_o�_�_o!o3o Uo�oio�o�o�o?_�o �o�o	7?mS e�����oZ�Q �Vy�Wy