��   ?Q�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����MN_MCR_�TABLE  � � $MAC�RO_NAME �%$PROG�@EPT_IND�EX  $O�PEN_IDaA�SSIGN_TY�PD  qk$�MON_NO}PREV_SUBy �a $USER_�WORK���_L� MS�*RTN�  %SOP�_T  � {$�EMGO�}�RESET��MOT|�HOL�l��12�S�TAR PDI8�G9GAGBGC��TPDS�RE�L�&U� �� �EST��^�SFSP�C����C�C�NB���S)*$8*$3�%)4%)5%)6%)7�%)S�PNSTR�z�"D�  �$$�CLr   �S���!����� VERSION�(�  ����!IRTUAL��/�!;LDUIM�T  ��� ����4MAXDR)I� ��5
4.�1 �% � d% ��}? i?�?���" ���?�?�? O�?�?6O �?3OlOO-O�OQO�O uO�O�O_�O2_�O�O h__�_;_M_�_�_�_ �_�_�_.o�_Rooo Mo�oIo�omoo�o�o *�o`�3 E�i����&� �J�������}��� e�w�쏛����я� X�C�|�+�=���a�֟ ����џ�͟B��� x�'�����]���䯓� ���ɯ>��;�t�#� 5���Y�ο}����� �:����p�ϔ�C� UϏ����� ߯���6� ��Z�	��Uߢ�Q��� u߇��߫� �2���� h���;�M���q�� ����.���R��� ��������m������ ����`K�3 E�i����& �J��/�� e���/��F/ �C/|/+/=/�/a/�/ �/�/??	?B?�/? x?'?�?K?]?�?�?�? O�?�?>O�?bOO#O ]O�OYO�O}O�O_�O (_:_�O#_p__�_C_ U_�_y_�_ o�_�_6o �_Zo	oo�o�o�o�o uo�o�o�o �o�o hS�;M�q� ���.��R��� ��7�����m���􏣏 �ǏُN���K���3� E���i�ޟ�����&� �J������/���S� e����ׯ���ѯF� ��j��+�e���a�ֿ ����ϻ�0�B��+� x�'Ϝ�K�]��ρ��� ߷���>���b��#� �ߪߕ���}ߏ��� (�����#�p�[��C� U���y�������6� ��Z�	����?����� u������� ����V S�;M�q� ��.R �7�[m��� /��N/�r/!/3/ m/�/i/�/�/�/?�/ 8?J?�/3?�?/?�?S? e?�?�?�?O�?�?FO �?jOO+O�O�O�O�O �O�O_�O0_�O�O+_ x_c_�_K_]_�_�_�_ �_�_�_>o�_boo#o �oGo�o�o}o�o�o (�o�o^[�C U�y���$�6� !�Z�	����?���c� u������ �Ϗ�V� �z�)�;�u�q�� �����˟@�R��;� ��7���[�m�⯑�߯ �ǯٯN���r�!�3� ������޿�����ÿ 8����3π�kϤ�S� e��ω��ϭϿ���F����j��+�
Send Events��S�SENDEV�NT��Q����� %	��Data<�߶�DATA������%��Sys�Var;��SYS�Vw��ڗO�%G�et�x�GET�+��%Re�quest Me�nu���REQM'ENU?��ۚ�]� ��Y���}�+����� .��d�7I �m����*� N�����i {��/��/\/ G/�///A/�/e/�/�/ �/�/"?�/F?�/?|? +?�?�?a?�?�?�?O �?�?BO�??OxO'O9O �O]O�O�O�O___ >_�O�Ot_#_�_G_Y_ �_�_�_o�_�_:o�_ ^oooYo�oUo�oyo �o �o$6�ol �?Q�u�� ��2��V����� ����q�������� ˏݏ�d�O���7�I� ��m�⟑���ݟ*�ٟ N������3�����i� ��𯟯�ïկJ��� G���/�A���e�ڿ�� ���"��F����|� +Ϡ�O�aϛ������ ����B���f��'�a���]��߁ߓ��$M�ACRO_MAX�X�������Ж�SOPE�NBL ���2��ݐѐ�_����"�PDIMSK��2�<�w�SU����TPDSBEOX  K��U)�2�����-�