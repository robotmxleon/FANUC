��   ��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����BIN_CFG�_TX 	$E�NTRIES  $Q0FP?UNG1F1O2F�2OPz ?CNE�TG  �DHC�P_CTRL. � 0 7 AB�LE? $IPU�S�RETRAT��$SETHOsST��NSS*� 8�D�FA�CE_NUM? �$DBG_LEV�EL�OM_NAmM� !� FT�� @� LOG�_8	,CMO>�$DNLD_FI�LTER�SUB�DIRCAPC � D��8 . �4� H{ADD�RTYP�H NGGTH���z �+LSq D �$ROBOTI<G �PEER�� �MASK�MRUv~OMGDEV�����RCM+� 7$ �/�QSIZ�T�IMR� TATU�S_/!?MAIL�SERV $P�LAN� <$L�IN<$CLU���<$TO�P7$CCw&FRw&Y�JECZ!8%EN�B � ALAR!B�TP,�#,�V8 S��$VA5R�)M�ON�&��޶&APPL�&PAp� �%��'POR��7#_�!�"ALER�Tw&G2URL �}83ATTAC��_0ERR_THRO33USt9&!u8�� CH- A%�4MA�X?WS_Z1���1MOD��1IF� $�2M (�1�PWD  } LAطr0�ND�1TR=Y�6DELAC�0<%'�1ERSI��1v/'RO ICLK=HqM� /'� XML+ ��#SGFRM33T� /!OU33PIN3G_�COP�!�F�3�A/'DUMMY�1�G2��RDM�*� $DIS��SM !l5�M!n"%/7�I�CC�%� FVR�e0GUP� _DLVNSPAR�QN�
#	3 _)R/!_�WI�CTZ_INsDE�3�POFF� ~UR�YD��Sk � 
 t �8!]PMON� cD\�bHOU3#EA�f.af.a%fLOC�A� A#$N10H�_HE���@I��/ 3 $ARyP&&�_IPF�#W_ O�F�PQ�FAQD0�VHO�_� INFOncEL� P����0WOR�1�$ACCE� LV�5[02�ICEد'p �$�c  � Fq��
��
�;p&PS�ADw�# ��WqIX0A�LCUq' dx
�
��F����op�r�uw�$� 2�{���Qr�}�p�� ğ}��!Mq5����$�� _FLTR  \cy�p ���������I�$�}2�I��bSHyPD 1}�y  P1�珴t֏��7��� [���B���f���ٟ ������!��E��i� ,�>���b�ï��篪� �ί�A��e�(��� L���p����ҿ�ʿ +��O��[�6τϩ� l��ϐ��ϴ����9� ���o�2ߓ�V߷�z� �ߞ߰����5���Y� �}�@�v���������M�z _L3A1�b�x!1.6�0����5�1F���2�55.~�=�����u4�2;�M���a�s�������3��M�* ��������4+M��  Qcu���5�M�@������6�M��ASew����$RC�`G �MA� MA���Ѐ�v� OQ� ���<-/ b/t/G/�/�/�/�/�/�/��P�/"?4?F?? j?|?�?�?_?�?�?�?��?��u2OLO��?wO�O�O�O��}�iRConnec�t: irc�D//alerts�O �O__*_�EqOV_h_�z_�_�_�_���sP�"��d���_�_�_ o!o3oEoWoio{o�o�o�o�o��$E_�o��(�oiO:L^pR����(�$"��r&J�u�q��� D�M���$SM&��ŋ��%1�D���I���8�q��\��� L�qN�q
!	��~��珿�p������ #��US?TOM 
�}����#  ���T�CPIP�r�}�$H%�TEL���u !� �H!T��R����rj3/_tpd�� $�ׁ?!KCL�����׏��v!CRT����W�"ߔ!OCONSX���őOsmon]�ߔ