��  U��A��*SYST�EM*��V9.0�055 1/3�1/2017 �A0  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ���AIO_CNV�w l� RAC��LO�MOD_T�YP@FIR�H�AL�>#IN_O�U�FAC� gINTERCEPf�BI�IZ@!LRM_RECO"w  � ALM�"�ENB���&ONܢ!� MDG/ �0 $DEBUCG1A�"d�$3A�O� ."��!_IF�� P $E/NABL@C#� �P dC#U5K�!M�A�B �"�
� O�G�f d��APCOUPLE, �  $�!PP=_D0CES0�!e8�1�!��R1> Q�� � $SOF�T�T_IDq2TOTAL_EQ� 3$�0�0NO�2U �SPI_INDE�]�5Xq2SCRE�EN_NAM� �e2SIGN�0�e?w;�0PK_FI�0	$THK�Y#GPANE�4 �� DUMMY1"dJD�!UE4RA��RG1R� � _$TIT1d  ��� �Dd�D� �Di@��D5�F6�F7�F8
�F9�G0�G�GPA�E�GhA�E�G1�G �F��G1�G2�B!SB�N_CF�!	 	8� !J� ; 
2L �A_CMNT�?$FLAGS]��CHE"� � EL�LSETUP �
� $HOMEm_ PR<0%�S�MACRO�RREPR�XD0D+�0���R{�T UTOB� U�0 }9DEVIC�CTI�0�� �013�`B�Se#VAL��#ISP_UNI�U`_DODf7{iFR_F�0K%D13���1c�C_WAxqda�jOFF_U0]N�DEL�hLF0pEaA�a7b??a��`$C?��PA#E�C#sATB�d�� oW_PL�0CH/7 <� PU�P��B
2ds�`QgdsD�UT�PHAgpS�F���WELD|H2/0 =Lc�7w7atAING�0�$�r�1�@D2�4%$�AS_LIN;tE��w�t_��2UCC�_AS
BFAIL��DSB"�FAL�0�AB�0�NR�DY��P�z$�YaN�Wq<��`DE6r ��`���+�����tSTK��+�;s7�;sNO�p��[�̈́r��U* Ȁ%�9 � ��  ��q`�G�C�G�+�U�S_FT�vpF�ǂG��SSF��PAUS����ON7xǓHO5U�ŕMI�0�0�ƔSEC�2�ry�i �rHEK0�v8vG#AP�+�	�I� � gGTH���D_I���T= �l���� �`�s9!̅����9!G��UN1���q���#MyO� �cE � �[M�c����RE�V�B7��!XI�� �R  �� OD�P-��dPM� %�;�/�"8�� F�q��
aX�0DfT p{ E RD_E%�~Iq$FSSB�&_$CHKB�pEde#AG� �p�  "
�$Ա� Vt:5���3�Mpa_EDu �� � C2��qS��`�vl �d$OP��0�2�a<�_OK<��Y�TP_C� <�pd�vU �PLAC��^}��p� xaCOM	M� �rD|ƒ��0�`��KO]B BIGA�LLOW� (tK�w�0VAR��xd!�1}!�BL�0S � ,K|a�r�PS�`�0M_O]|=՗�CCG�`=N�! �� ��_I_��� �0�� �B.��1S� ~�CC'BDD�!��I����0�@��84_ CCWp` OOL
��P'�M�M
�n�CHs$MEAdP�d`T�P�!���TRQ�a�CN���FS3��ir�!/0_F��( D�!��v CFfT X0�GRV0��MCqNGFLI���0UJ�p����!� SWIl��&"D�N�P�d��pM~� � �0EED��!��wPo��`�PJedV
�&$�p��1``�P��ELBOF� �=��=�p/0���3P�� ���cẐ�G� �>A0WARNM�`ju���wP��𼠤 CO�R-�8`FLTR^juTRAT Tlp�� $ACC�rT�B� ��r$OR1I�.&��RT�P�p\gMpCHG@I��E3�T{�1�I ̉ra�HK��� �����"�Q���HD(���a�2
BJ{PCT��3�4�5�U6�7�8�9�!����COfS�_rt���3�V�O�LLEC��"MULTI�b
2��A�
1c�O�0T_�R � 4� STY(2�R���).��pp�b�n� |A0@6Kb�Ib$���P�c���UTO=�cE�EXT!Y�
B�!�Q 2 
l��a0��Rpub����  �" ���Q����qc��~#!|��1Y�M�
�P8$  lT}R�� " Lqࠊ/��P��`AX$GJOB׍��W�';IGx# d��? %?78��3�p%���9_MOR��$ et��FN�
CNG&AF�TBA���6䱀JC��9��D@r��1CUR.KPa`/Ek��%��?��ttaoA4��XbJ��_R��|rEC�LJ�r�H�LJ��DA���I�����2G���]QCRfT&�C ��bG����HANC6$LG��iqda��N�*�Ya�Cᇁ�0|rf�R'L±�mTX���nSDB�WnSRA�SnSAZ��P�X��$  ' FCYT��e�_F��Pn�Re�M
P�QIkOh ������1��e����Cg���A���MP�a� ��HK�&AE�Up�p�Q�QI�'�  ]PI���CSXC��Zq( �xs��s��T�R�C�cPN����MG�IsGH"��aWIDR��$VT�P��9�E�F�PA cI�X�P,aQ�1u�CUS�T��U��)R"TI�T����%nAIOV����P_�L����* \q���OR��$!�q���-��OeP��jЅpIp�Q�u��J8�
��0�_�~}pPXWORK��=+�$SK0���nWADBT)PTRw�_ , �l@Ab��s�R0�ؠD��A:0�_C����=�+`H�PL�q��R�A�"��#�D��r�����BJ�b��9�����DB�Q2��-�r~qPR��ΰ�
x ct��. p�E�S�a� �LӉI/��-�( ��0���j� 1%��EsNE���� 2D��b��q	����3H�PC�  .$L��/$Ӄ�����gINE׶�q_D����ROS��E0"2`q��f0�p��PAZ�|tAsbETURN�����MRQ2UA@�C�RŐEWMwp��S�IGN�A&rlPA���W�`0$P�f1$P�P� 	2j���q����!��DQ��f������׶GO_AW;0���pvp��qajDCS'����CYx42O�1P�8�8���2��2��N�@��CtDۣDE�VIѐ 5 P7 $RBֳ���I�P.�i�I_B�Y�q���T�A9�H7NDG�6���x����b�DSBLr3�ͳ��aܢLe7 H �� ���TOFB̶�FE@Бg')��ۣ�f8��cDO�a�� MC9�@�"�`�sr�(��H�P�Wp�X�ܢSLAt4���9IINP!���� ж�ۡ�:D *�SPNp�#�@lƍ�1��W�I1��@J��E�q87�qW�N�NTV#��V n��SKI�STE^�`�b��pڥ�aJ_�Srjb_>���SAF��k���_SVBEX�CLU��po�D�pLX ��YH��%qΉ�I_V9`�bPPLYj���������_ML��L�VR�FY_D��M�IO�`  P�%`�b�Oe��LS�|b��%4}������aP�u���Y�AU NFzf�����)��#"�cD�4Ͱ� S��r�AF� CPX٣e�_� ;j��pTqA#���  ��SGN��<��<@3� P��c_�t�a���qd��rt��`UN>�����<@rD�p]�T`��`��%`����zrEF�p]I>�= @��F��\t6@OTS����|�������孂y Mr�N�IC>2K�GM A���iDAY�sLOCAD���D��5��o�EF pXI�%?j���~cO� �5�_RTRQU�@� D����0Q�p �EԠ��� �?K�%>`� ��GAMP*Pp��A�"�'; DB'��VDUtS�U��CABU�B`�NS9@ID�1WR$�Q!`�V[�V_#� ; ��DI@J$C� �/$VS�SE�#T �BDC�A� ���|�DBf�AE_�;VE�P�0SW!�!�@�x�3�� @�`�O�H�@PP <I	RwqDBB�p�=�!pU����t"BAS�рo'~P�Pn%[�d� B�	� ���RQDWf]%MS� �%AXC'<�;LIFEC���� ��	2N1EB5��D3EBCd@/Ź�Cq`ʡN�4q�6��3OVՐ%6HEh�DB'SUP�1��	2D�_�4j�H1_!C�5š
�7Z�:W�:qa�7�S��"BXZ�PʁEA+Y2HC��T�pސ��NM��zr0P�dgD `L��@HE�VXCSIZ?6k0��[��Nh�UFFI�0���C��������6ܭ�HMSWJEE �8��KEYIMAG�TM���S�A5���F���r��OCVI9E �qF 	�P�LQ�_��?� 	��&`KDG� ��ST��!>R|�FT���FT� FT� FPEMA�ILb �aA|p�FAULSHR�*��;pCOU_��q|pT���U�I< $d�S_�S#�ITճBUFkG�kG@�jpJ`p�0B�Tk�C�p�Rws�PSAV(e �R�+Bd�$ Cg�p��AP/d_ň�$̰_�Pec �iOT�����P@����jA�gAX��sq:p�P��\c_G:3
�YN_e!�pEJ0Df�W�r�d"UMO_0T��F�� �E2���^Јq	K��ey&^�5rH 8)�4��qL���nqL�S�cC_ܐ��K��pu�t��R�A�u�X�nqDSP�FnrPC�{IM5c�s�q�nq��U�w{0�0��PI�PR�nsN!D�@�sT!H��"ûr� Tߑ�s�HSDI�vABSC_�9@`�V��x�v���c~����NV��G ��~�*@�v�PF!�`ad�s0p�a��SC��\��sMER��nqF�BCMP��mpET��⌐M�BFU�0D�U�P?�M�B
�CD�yH��`�S9pR_N)O�ዑN� %�i�Xcg��PSf�C�@%v�C���a~Qd��`U OH����c  d�������}�锍� �9疗疢疮A*�7�8�9�0T��1��1
�1�U1$�11�1>�1K��1X�2f�2���2�
�2�2$�21�2�>�2K�2X�3f�3R�3��
�3�3$�U31�3>�3K�3X�94f��QEXT�TP <sK�p<6p��p2ǋ��QFDR^�QT�PV���b	2p�v�	2REMr�F��0BOVM�sz��A��TROV�ɳDT3`��MX��I�N��Q0�ʶIND����
	�i��`$DG�a{#��4P5�9D���RIV"�=2�0BGEAR�qIO�K��;N0p}ة��(���@�0<Z_MsCM@	1 �F|0;UR"�R ,t� a�? P0�?\��!?��EG ��`a��e�SG � 5P�a�RIM��@��SETUP2_ gT � �STD6� ��<����I�C�`��RwBACrU T[ �RTt)Nz%��+p�IFIQ!+p��А���PT{b[�LU�I1TV � Y�PUR�!�W2�r�<qv��P�� I��$��S��?x#�J�QpCOw`�cVRT|� x$SHO���SASSY��a?5P8�W����A�W�RKFU��15q��25q���*@�X |�N;AV�`��3����*@�R=1��VIS�IJД�SC���EP�c�\�AV��O���B%EX�$PO��I\ ��FMR2b�Y o�X�}p� bpNt�{ߍߟ߶ơP����_f�G�_���B��M4�Y�k�D�GCLFR%DGDMYLD��7�5!6H.�04%�MR�3SZ�@��	 T�FS�`2T[ P!��bs>�`$EX_��B�1�`Ā\2�3�M5��G��9\��
���PWeO�&D�EBUG��"��G�RR�spU�BKUv�O1�� 0PO� ;)' ��' �Mb�LOO�ci!S�M� E7b������� _E ] ��@Y� �TER�M�%^�%[�ORI�Bq� _�%1SM_OpL� `�%^���(�a�&�@UPRbg� -���]�#0^��G:0E�LTO{Q$US]E��NFIc1G2���!���$4_$U;FR��$j�A1�}0=�� OT�7��TqAX�p��3NSTCp�PATM�d@�2PTHJ�;�E4P_bD�H2ARTP`R5�PPa�{RG1REL�:�aS�HFT?�H1�1�8_�N�R�8��& � $�'H@a�q�B���b�SHI@�U�� JaAYLO��a�a����Y�1��~�J�ERVA�3H7�Cp�2�����E����RyC�~�ASYM.q�~�H1WJ[7��E ��1Y�>�U2TCp �a�5�Q=��5P��@���bFORCpMKT�z!:c��'"`&0�0w0�a� HOb�f�d Ԟ2��& X�O�CA1E!��$�OP����V�t �����P��P��`R�Ń�aOUx��3e���R�5Ie h�1��eo$PWRL�IM;e�BR_�S�4��� �36H1UD�_C�RBt]e7�$HSu!�`�ADDR2�H}!G �2�a�a�a��R��x�f H!�S����u��u
�u�SExv���!�HSH��:g $���P_�D�H Y�RrPRM�_��^HTTPu_i�Hx�h (*��OBJ���b��$�2�LE�3�s�i� � #�"�AB%_
�Tp#�rS�Px����KRL{iHITWCOUw�B6�L `�rQ��U�`��`�SS��JQUE?RY_FLAQ1�pQWR�N1x�jpgP&��PU����O���q��!t��/t����_�IOLNw�k(��� CJq$SL�L$INPUTM_Y$;`��P,���C̀SLA� l׀�(�$��C����B1IOgpF_�AShm}�$L ��w��8AِU� 4@�_1��݃��情@HY�1ǧ����a[�UOPen `l�ő2��� �������[`P�c;`��	������NqUJ�a�o � K�N!EaG4�v7F�Da��2�J7VpOQR$J8q�7�I_1z���7_LAB�1�P|����p�APHI���Q{���D�J7Jx�-��_KEY�� �K��LM�ONx�p�$X�R_���)�WATC�H_��C��D�EL�D��y����eq �@Р1V�@&�U�CT�R�3U�i��*l��LG��r� !#�LG�Z�Rࢵ�c��c���FD��I ����\!����� ���� e�Dqf�ce�c�e�ΰ�e�� e���@0J_@�ѐ1j��qʦ�F�A�xǒĞ�Cd(��SB����c��c���ΰ��I�����ƍ ̷ƞ�RS��0  �(ʀLNe�<sѐ���)��6�"��UosD��PLM�C�7DAUi�EAwp���T�u�GH�R1o��BOOw�t� C���`IT\���� 8������SCR���㖇�DI��Sw0HRGX ���z�d(��o���w�W�o�X��z�JGM^�MNC�Hl�n�FN�a�Kn��PRG��UF���B��FWD��HL.��STP��V�� X��Г�RS�HzP��w�CdD��1Rz�: :�^�Unq��9���H�k�����Gw�@( w�`������s�}�OC/ v��EXv�TUI��	I��7�C�O������<@���	$���<@��NOANqAo�A2� VAI����tCLUDCS�_HI$�!s�O��
�SI��S��IGN���ɳ��h�Tc�DEV�<�LL�A��_SBUI �uP�j@mT��$��EMr����]���*"	1vP�@j@ހ��~p����1�2�3�>��� 
0w �C��x�Q@5������IDXa$9 [�����֥1�STƐR��Y� <@   v$E.&C.+�pmp�=&P&����	1x L ����`��4@r�`Na��eENwp�dp��_ y ap7�}px	b���# �MC7��z �C�CLD�PƐUTRQLI��TT�94FLG )"0�Q53�DD�57�t�LD55455ORGT�8�H2_ȲF�8!s�D/r�#�S{ �� 	59�455S�PT0��0y0�4}�6RCLMCD@�?�?Iƀ�1pM�p�^���|�$DE�BUGGugQDAT�AY��T �UF�E��T)!��MI�6p�T} d@��R�Q��0DSTB��`� �F��HA�XR��G�LEXC#ES$R>��BMZ`��~� �B4���BSq*�����F_z@�H��S[�O�H�MJ;PTH�� &Pv��m��QMIR� �s � []R�WRCT��N}��VUO�ZA�ZL�RC�PQC��Q�`D��O��^�CURPX_THqG�P�`R`|1�o)`/d55R^`�`S<�P �B_FR@^�a\fZ_��^ddpG���* �!KH�� \���r�Fv$MBu�L�I�q�cREQUI[REG�MO�lO�k�fB�$ML� MG�� ap���`|��cB��ANDU�Sz��>�5�Z�9sD��Q�IqN�p��Q�RSMf�(Sx� �Q�!E]�q�RA'qPST� 7� 4�LO�P��RI ��EX�vA�NG��AQODA5QG���@$�QG��MFh������"���%&�2ТfSUP��%4QF `RIGG>�� � ��0�#�1��Ӫ#Q��$$���% #n�א~�א��rP��8wAZw@ETI9�~��Q2�M\p9� tV�pMD�I��)��� �DA�H�pu���DIA���ANSAW,��w���D���)�!O7��0�Љ �QU��VB�70�B�L�p�_V@�ъ ��C���sX@�b|�ٰ��P���v���Pƴ�KES�!���-$qB����� ND2FB���2_TX�$XGTRA�1����`LO�ЪЋ$RG��B�F�8Ҍ|�g�_��4RRR2�E�0� #W�e�A�1 ?d$CALI�@2��G���2�RINܩ���<$R��SWq0"DᣫABC�x�D_J��a����_�J3�
�1SPHs�P��P�-�3,�(��?���\�J�l�4�2�1O8IM� �2CSKP":��~�Y���J���2Q��̵��8̵·�p_AZ�2h����ELg�FAOC�MP�s�1!I�RT�A)�Y�1�i�G���1�K�> Y�ZW�ScMG�܀�4JG� �SCLP�uSPH�_� �0����������RTERࠧ�o�IN��ACz��|��� ��r��} _�N�я������2L4��?R� �DI�OA��DHP3��ё�$V��Rs��>$v��p�1�����@Ro��ВH? �$BEL�?w~��_ACCEL�a�ث���P_RـJ� �QT!�*aEX2L6b��3�� �׀c��.a�����-36cRO
Q_�m��J�P��2�p`��_M=G�$DDm�����$FW�0݀�Ӱ��Ӥ�~�DE��PoPABN��RO��EE`���0±�PYAOP��oa_��JYPaPC��YY����1 �!YN�@A ��7����7�M�A���ig�OL�de�INCa��q����B�����AENCS��Á�B��Ѥ��D+`IN"I�6b��ހ��NTVExk���23_U������LOWL�`#F�0��DF�D �`��� ��`RC����MOS� wT�PP�2���3PERCH  8OO`�� z�q� !�4!$��!�)b��A6b�L�tW�����F�
4TRK��!AY[�(cOQ I�XM�p/�SQ�� MOMc��BOR�0���D�㣧d���捠DU��7bS_BCKLSH_C� ��@YO`?�����*N�ĵCLALM����1�?P6%CHK�0� �GLRTY@������Ѕ|1܁_�NN_UMzC�&CzCp{���#��LMT)��_L�0ú$+��'E �-� �+� ���%��>�0�C�!4�PC��!HI��`q�%C@8�\{��CN_��N"CL�6��SF�ѯ	V!�p!����U1��5Y8CAT�.SH���� ��?a���X�7aX�L�fn�PA�$��_P�%s_����Pn ��`�rDc%JAaPfC	 O�Gs7�TORQU �A�Li���bd����B_W�IU�nѠ�D_��Ee��EI�KI
[Ie�F�P�As�JX,��w�VC��0��jS1q^o��_��wVJ�RKq\�R�VDBґ�M��MPp_D9L_��GRV�D�T0_��Te��QH_^��S�#jCOS0k1�0hLN�PSktUZd_�Ui�v�Ui'Q�jlEQ�UZN`d�QMY\a�h<b���Dk�iTHET0$NK23e�rYӶ]`CBvCBY�C��ASrqDr'TRq_ӌRqvSB_�pr*uGTSֱ��C0��qO��;C_Ǧz�c$DU ` ��r����xR�v��b�Q��53�NE��7�I^`q#;��=�q�Au;�D�"e-h-aLCPH0e����StU ��e���e��f�����f=�V]�VR�O�u�UV��V��V��V��UV��VɋV׉H]�@��|�t��1����H��UH��H��HɋH׉�ON�O]�O�s�O���O��O��O��O*��OɋO�fF�?q�e��P�SPBA�LANCEc�=1LmE�pH_uSP���pf�f�fPFULC������e��{1�+�UTO_[ ��ET1T2_���2NB!�����у �P�p�ҚӞT
O�|���@INSEG�Ҏ=REV��= ��D3IF3�1��1�1�&OB�&!�S°2�@��M!�TLC�HWAR��T�AB�BA�$MECH`Hq�`V�\�q&AXV�P4u�4�@�T�� �
v��Ab���ROB�n CR���j2?�MSK_֠��_� P j�_�AR���2����51�2���������$��>�I�Nű�MTCO�M_C\P�Д � h���$N'ORE��Q��.�@�o� 4�@GR�B�a�FLAű$XYZ_DAQ����/DEBU���f�.��mЖ �$/�COD! �҇b���$BUFIwNDX��  ���MOR��� H �����E&��~�^�$޲��o1�� CTA�����ҰG���� � $SIMULp@�С��\��OBJE��\�A�DJUSz�m�AY�_I�A�D��OU�T�@�Ԡ_�_FIb�=��T�@���� ����q��������:�D,�FRI��MT�RO�@��E�A>�OPWO�P����,��SYSByU+���$SOPT����;!_�U^��PR�UN0҅�PA��D��`�Y� _��2z���AB��
0��IMKAG!���Pϱ3IM���IN�P��~��RGOVRD�v�e��P����� ���L_R�zA(�"�0R�B� � 1MC_SED��b� 
0N+��MW	1�MY19n1��SL������ ���OVS�L��SDI5�DEAX�3��3
�V�@�N��A��� ��(�n�C�0T�x�6�_SET�@��� @�@!��CRI^���7_Lq�@YLc��x�0 ����Ta��@AT�US�$TRCp���ҔBTM��I��l41sU .��� D��E���4�E���� & �EXE�r!L�� "�)�0���U�P��!IS��X�NN��1ldQ� ��PG>՟L�$SUB��V�Z�JMPWAI�0P��%LO� ��̰[��$RCVFAIGL_C�i�!R�� i�r�e1�0�4���%�`�R_PLZDBTqB�A�2i�BWD�&fY�UM�@�$IG��8�����0TNL�0�$@2R'�T�~@�@��P�PEED5 �3HA�DOW�@c�Y�f�E��4�p!DEFS}P�� � L���|��0_�0���3UN!I����0C!R iL�`̰P���	P1�����Ю@^Ѻ��� ���N�KEQTB�@��	@P42���� h �pSIZE��������`A�Sx�ORZFORgMATK�*4CO~ ,\AǲEMn�|D�3�UXC��p�PL�I%2��� $I�O?MP_SWI/��%E��Wi�JscѺP�
0%0AL_ ���@�0"�gPBJDpC��D��$E!��J3D�H� TV@PDCKC m�CO_J3r�RQR�Ģ�	_]��@C�_/1A  � ��h�PAY�qҧT_e1�Z2�S�@J3�p��[�U�V�S6�TIA�4�Y5�Y6�MOM�c$cc$cc;�B� ADcHfcHf6cPUSpNR)due�cuebm"�A�ħ?` I$PI��U lq�U*s�Uus�Ujs�U Ut�f�kit�t��v��v_!��m����v3HIG�Cv3�%�4iv �4�%� ��iv�sxx�!8�y�!�%SAM���p�tiw�s�%MOV��$�'�
�ް)p%�� � #��0�P2��P%�0� 5�`!��@��H��#�INj��@�sq���h���"s�������ӋGA�MMǦ���$G#ET���Є�D�T/�=
z�LIBR9!W2]I��$HI8 _��H�%�H�E"�U�AO�r�c�LWJ�����r�@��c��Rn�M0�AC5x0� a ?^I_�p2�/��B�X�A�Y��$c/�Hf��C ��$,X 1U���IXRk�D�0>�A!�$@�LE �8q�`���Xq��Z0MS�WFL�$M�@SCRI(7���)q�T"p�0�A����P���UR�$�v�KS_?SAVE_D-B�;#NO�PC`<"�T B�&��_�a�YW��i�Y �`����pkR#uܸ�SD��p#�s0�@�,� $�cxY�sv�x@�<Š���<!>��@M�ũo � "�YL�c��Y��S��6�0 �� 0����J�������H�	�t�Wq�����`��1�t�M����CAL���Q��o �1T"�@M3�*� � s$��G$WR� �����QR�oTP�vT P�}TP�T0���+�(�C;�@X�0O~S�A�Z�տ@��Uԫ �ՑOMK��V����p����̿`CON��� �c�Q_v"� | =Q�B�$i��c��c B��Z���j�A �x�(������P���P_A�PM� QU��p � 8@Q�COUM�i�QTH�/0HO��G�HYSf�@ES�F�UE2�t8�E@O�D�  �@1P0�@�`UN������OVr�а P�����%$��W2RO�GRA���2�O�����IT����t�IwNFOXѱ �A8��������� ((�SLEQ�Zv/Nu/ ��N�OS���s$� 4@E�NAB~�� PTIONZ�4(r��4cWGCFl�0J� ��A���,�R��� +S_E9D� �е �N�ЩK�[sG�E��N9UAUT^�COPY�8 7�1�j�MN�NAE�PWRUTf� HN� �OU�B�0RGAkDJXѶTBX_t���2$�0��мW�P����v3��#�EX� YC~��-
�NSh���ޠ�LGO��PNYQ__FREQ�bW��0MvM!�D��LA��D!p�c��[uCRE3��R���IF�a��NA��q%�$_G}4T�ATB0�$>�MAIL�r2��!��B��1�!�1�$ELEMl�� �s0vFEASIy@���@��2[q K�66�V�2�I��0��D"8qJ��k2AB$�APE��vpV�!�6�BAS&R�52��aU8�p��W�$�1�7?RMS_TRe3�A����3�ӓp�r�!�4 �  !"�����	~B2 2� �� �ԇ�(F�2'G�2/�_�����2SG�g��DOUd��N�!"PRe�zm �6GRID���b�BARSZwTYHzp�U�O?`Xѻ�`���_�$!��B�DO|��i� � ����POR���C�f�B�SRV� )TVDI`�T�P0QCT� MWTCpMW4KY5KY6KY%7KY8/Q�F�l���$VALU��35�(42��Fh�� uY����C1�!2�� AN4��R�!RR!2�TOTcAL�s�a2cPW:#�I�AHdREGENFj[b��X�8��R%��V-�TR�3�rFa_!S8��g[`�V���b��2E�#�@L�1¸��-cV_H�@DqA-��`pS_Yf����^&S�AR-�2�� �IG_S!EC�`R�%_���d#C_�F�Q�E�q�O8G6�kjxSLGEpl�� >�_%��/�0`�9`S���$DE.QU0>���  �pTE���P�� !�a��a�J�v^�3IL_M`m$;����`��TQ-�6���0Ƨ��Vh�C�v�P�#1��M��V�1��V1��2��2���3��3��4��4 ��$��`ӓ%�� 0���v�INA�VIB=�Pp�]��d�2`�2l�U3`�3l�4`�4l��X�WB�qB����D $MC_FP���%�LC�B�f�#cMo�I��oC ���6��q��KE�EP_HNADD"�!#��0-�C�ѫ AC��A⒤�D�O&� "�{��3�D��!a#D�REM[�C�8a�B�������U�$eC�HPWD  #��SBMSK�BCOLLAB/��P@�$a�" IT$ ��f�ȕ��� ,(�FL�{�W�M�YNڐ1�M���C`r�G`UP_�DLYX���DE�LAc�9a�"Y�A�D-��QQSKI�Pw�� �P��OƠ�NT9�����P_ �����ҏ�÷�a ѹ�ѹdPкqPк~P�к�Pк�Pк�Pк9���J2R ���
qX�0TG#r���q�r�� �r����X�R�DCS�� �_�R"�R1�o�=�R�!��8J��*DRGE� T3�ÆBFLG'�����*DSPC��!UM�_r�!�2TH2N�rA<�e� 1�� 2��@� 11��� l����O�v�ATy��.��Q& �������� *D�Ҙ�B��H��ҥV�2]ҁ�c�u߇ߙ߽߫� +�U�3]������p��(�:� U�4]��]�o��������5]��������P�"�4���6]��W��i�{������� 
U�7]��������
\. NU�8]��Qcu������S�L�  @�1V�p`�L㙠E%$рp�e)fcIO��Ip���POWEC�� 1M0���N�#d� �+��$DSAB] � �""c^�CBД���M
E�+��	D���0E�"��MD8"' "�D� D�p�'/DBG_~@PD�3L%!eaPG
A@����@S232i֓ ����P��pI�CEU�2!`k$�pA�RITq!aOPB��rFLOW>pT�R(.b��@qCUz� M%3UXTA��qINTERFAiC�$��U`�v� CHA� t�0ݐ"!hp�$�`�`�OM'p�sA���0IHᓴ0Q@A+ӪTD�Sv`���8c3�E�FA����r�S�# k��`8b q��Rq H��6A ٶ��q  2� ��S��M �	� �	$)�s�0�
eC2`�_%pFDSP)FJcOG�`�#�p_P���"ONg�u���'�	6=Ky0_MIREAb$fwpMTY��CAPK� wp4Ц@�4"ASp}@�r"At �EBRKH <16=��R�� �B�s��BBPo0�bC@B�SOCF��NUD�1pY16��$S}Vi�DE_OPGt�FSPD_OVR��k��DTRWCOIRbW� N�PcVF�@l�WB@OVEESF�Z�^p�S,rF�V t'�U�FRA�ZTO�$LcCHa�u�2�OVST��B@WQ���BCZ� rx&PQ@]s  @��TIN�``!$O�FSC`C�0@�WD�|QdxQ%Q��E?PTeR�!e"�AFD����AMB_C��bB5@B<��!q�b�a�cSV��L�k0��s��R�G�g�HAMtB_0=0�e-b_M�`2x�:`T$CA8@��D�B?pHBKXo1~6TqIO�cu�pqPPAWz�qhy��t{uu�:bDVC_W R#�p1��p��@�Q�u���x-s�u3�v@3`��{�0p@SQUR#7@~CAB���,Ӡ�`���`�h9�O�`U�X~6SUBCPU�O@S������dp0�ݱ���c�d���$HW_C]��0ݱrp�ʆ�� �Ð�$�U��D���AT�TRI�0��O@CY{CLw�NECA)���CFLTR_2_�FI�/���L�P[KCHKՠ_S�CT�CF_�F_�|��FS��b�CHA��d����b�"��RSDU��Q�3��_T�hY���c�� EM"��M�CT���ݰĀ����2�D�IAG5RAIL�AC�sx�M��LO�	P7�/V���3� XH�3��sPR�pS+Г 90��C�q� 	^,cFUNC��1'RIN���$D���L�!ʰS_"@*?p�䣸�Mt���MtCBLȰ���A�
��
�DA�@�O���LD`0GPpqw�*A�|�w�TI����A�Ā$CE_RIYA��AF��Pn#Xò%`ȵT2d�C}3��r�aOI�fDF�_LY�Rl1�0LM�`#FA  HRDYYO�AM`RG|�Hސ�Q� W��MULS�E��3��8P�$�J_ZJzR�W�[FAN_ALMLV�#��WRN��HAR�D�@o6��2$SHADOW `I��@���V���!�Q�E_`�s�AU��R��2TO_SBR��6@�(�逺sá@�MPINF8`��S�m�^�gREG���DGy��K�Vm0��FDAL�_N�dFLۅ9�$Mm�l�J�g O`L��K$$Y�("V1�2#�o� ��CEG[�CGP
�A ~/U2p8S�;��EAXE,GwROB)JRED)F�WR  �A_i�SS�Y�@D��@��S��WcRI  �ɀST�P*C0�@nPE�&�w� �"@B��9a��5k�pOTOn�%`ARY)C�e����[@FI�@pC�$LINK�GT5H2��0T_��9a�%�69R[�XYZto2e�7s�OFFA``2� \�N�uOB'@�����a� h0��F�I���0�?T��AD_J�!�2lR?�pq������89R� ��	dT�AC��FDUWb�$�9x�TUR��X��z!�N�X��� )FL[��PH��� |����309ROa 1��KN@Ms�/U3���{�������W3ORQ�6A����{��@O��N��H�34A��N]OVEd("M00 J��~��~��}F1`|J�|�{AN�� 5�~ȱ)!e}@�� �ve�%��%��6AERSA�	|�E� �`��E$A�Ā���ܥ��V�S�V�AXc�2V��ҁ4�% 8��)b��)w��*�* r�*��*: �*q �*1� �&��)��)� �)��)��)��)��9�9�'9D189D7EBU��$����00��1VbV�ABV�Tq�|Q^VIp�� 
 B�s��+E��7G8Q7G w�7G�7Gr�7G��7G :7GqδF Ȳ4��LAB��)���sGGROB�)��2pB_�,&��uS��%���FQ*U�VAND� |�:$3�_�=!�YW 2qZ�^�mX�|X�5�^�NT��
c�PV�EL���QT��V��SERVE�P���� $���A�Q!�PPOHb���`��Q���R���� w $bTRQKґ
 ct�
`�gȲ2��e��Q�_ �� l���a��ERR���m"I� �P�raTOQ��LH�$�┅f�G�U%H�f� q  c��	a� ,�Q�#e=`��RA�a �2� d�b{s��S_a ����$r����"�eOC|G�p�  dk�COUNT�� �$�SFZN_wCFG	a� 4ƀ��;�T�Ŀ���3�����m!��PTq��� �(@M��o���`#������uFA���ö�sXd��{�y�aH��S��TO�d�PJ�?Y�SHEL��Yr�� 5k�B�_BASf�RSR�֤�^�S끐�M��1�gM�2p�3p�4�p�5p�6p�7p�8�g@�ROO��`9�f]�NL��LAB�S�N�N�ACKFIN2pTo���$U��M��� �_PUV���b�OU�P̠��-��f������&TPFWD�_KARwa��f`R�E�T,�P/�]��QUE���eU �����I��C-�[�[��Py�[�SEM3A�AA�H�A�qSTY�SOސ	�DI�ɠ}s����'��_TM��M�ANRQL�[�EN�DZ$KEYSWITCH^�s�.��ĔHEU BEATmM��PE�LEvb(��@��Ur�F�s��S3�DO_HOM�ưO���EFA PAR��rv����C���O8�c`�aOV_Mx����IOCMGd˗?�R.�HK��G� DX�׍pU��¹�M����HFO;RC��WAR(��b�.�OM� � Q@�4���U��P3�U1��2��3��4=�T rpO��L����b���UNLO9�����ED��  �SNPX_ASZr�� 0�ЄЍp���$SIZ��$V�AP�eMULTI�P��.�ŰA��?� � $H�/�H���B�S}s�Cr`���FRIFm"pS���������NFO�ODBU��~P������p�U�RN���� xU`SI�bTE�8��SGL*�TA� &�opC��C��+�STM�T�\�P��BW<e,�SHOWd�n ��SV7 _G�r� : $PC�@p7#֛!FB��P��SPbːA��� `VD��~�r�� �WaA00^T��ɰ��Ӱ���ݰ�����5��6���7��8��9��A��B�ٴ��׳A��y�B��F��70���1�U1"�1/�1<�1I�U1V�1c�1p�1}�U1��1��1��1��U1��2��2�2�U2"�2/�2<�2I�2V�9 ��p�2}�2���2��2��2��2���� `�>`"�3�/�3<�3I�3V�3�c�3p�3}�3��3���3��3��3��4�k	4�4�4"�4�/�4<�4I�4V�4�c�4p�4}�4��4���4��4��4��5�k	5�5�5"�5�/�5<�5I�5V�5�c�5p�5}�5��5���5��5��5��6�k	6�6�6"�6�/�6<�6I�6V�6�c�6p�6}�6��6���6��6��6��7�k	7�7�7"�7�/�7<�7I�7V�7�c�7p�7}�7��7*��7��7��7��*���P��Ub� Q`{@e�
n�V�ª�Q�U�PR��C)M�p�bM�PR9` ��TQ_+pR�P�e(a�~��SE�SYSL|�`�P� � L� �jw��A�ؠ; Ѡ�D��VALUju%�x���A6XF�AID_L���^UHIYZI��$FILE_L��Ti�c$��P�CSAq�� h �pV?E_BLCK���R|E��XD_CPU�Y�M��YA�us�_�T-�Y�*�F�R � � PW-p��<aLAj�SqAcRa�KdRUN_FLG de@dhaKdv�ke�a@d�aKeHF�Wd�`KduA�TBC2�u� � �Bk`(���ppĠ���d	�TDCk`�|r�b�p��
u�gT!H	�%s�D1vR��?ESERVE��Rt�	�Rt3���`�'p �X -$}qLEN���t	�}p)��RA���sLOW_��Ac1}qvT2�wMIO�Q�S���I.���B�Q�y�D}p�DE<���LACE,��C�CC��B��_MA�2��J� �J�TCVQ�r� �TX�s�����@����Ѷ� ���J+���Mۄ~�Jw����)�� ��q2��а�����JK(�V�K��:�>�:�sq/�J�0O�>�JJF�JJN�AAL>�t�F�t��n�4o�5/sX�N1�����d�N��DL�p_�Xќ��dCF6�� =`�PGROUDPFєQ���N�`C�� �R�EQUIR=rؠE�BU��yq܆$T��2�6�zp ��$�$CLAF� ����Z�*�*� qO���X�e����k�IRTU�ALW�i�AAVM_WRK 2 ��� ?0  �5a�ͯr٨ʯ�� ��A	s@�3�*����!�^�E�c�������`��ɿۿ㴧�BS�@��� 1x�� <��(�:�L� ^�pςϔϦϸ����� �� ��$�6�H�Z�l� ~ߐߢߴ��������� � �2�D�V�h�z�� �����������
�� .�@�R�d�v������� ��������*<8�~pN�LMTu�?���  dQI�NZlPPRE_EXE}� �~A�AT�ʖ���IOgCNVՒ~ �h�P�US���I�O_�  1��P $���I�4��1��?�?�`Tfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(��:�Q LARMRE?COV �c��LMDG �(BLM_IF m? ������+���N�`��r߄ߕ�, 
 �߾�9�E��������ANGTOL�  �
 	 �A   Y�k�Q P�PLICATIO�N ?�� ����ArcT�ool �� 
�V9.00P/0�3j�+�
883340����F0����1612�������7DC3��+���None+�F{RA+� 6��LP_ACTIV��	j��UT/OMOD� �Ո	�P_CHGAPO�NL�� ��OUPLED 1�  !3���CUREQ 1�  T=	=�=	�������=_ARC� Wel=�A�W�ՕAWTO;PK�HKY�D y�9'EK ]o������ 5/�/#/A/G/Y/k/ }/�/�/�/�/�/1?�/ ??=?C?U?g?y?�? �?�?�?�?-O�?	OO 9O?OQOcOuO�O�O�O �O�O)_�O__5_;_ M___q_�_�_�_�_�_ %o�_oo1o7oIo[o moo�o�o�o�o!�o �o-3EWi{ �������� )�/�A�S�e�w����� ���������%�+� =�O�a�s��������� �ߟ��!�'�9�K�`]�o����OTOC������DO_CLE�AN�����NM  H���^�p��������A_DSPDgRYR���HI��<�@M��&�8�J�\� nπϒϤ϶���������MAX��������
�X�������PLUGG�����
�PRC˰B:�"H����d�Oi�Կ��SEGF��� �� ����:�L��&�8�J�8\����LAP�� ��������������"�4�F�X�j�|�q�T�OTAL,�U�USWENU���� ߨ����O RGDIS�PMMC� ��C���@@M��O���߹RG_S�TRING 1~��
�M���S��
__ITwEM1i  n�� ������� '9K]o������I/�O SIGNAL�cTryou�t modej�Inp Simu�latednO�ut-,OVE�RR� = 10�0mIn cy�cl!%nPro?g Abor7#n�$status��${ cess F�ault�,Ale�r�$	Heart�bea�#�Hand Broke� ��/??%?7?I?[?m??��e��w �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O��O�O__�?WOR ��eKQ�?%_s_�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�o�nPOc�!�`c[ �o$6HZl~ ��������� �2�D�V�h��bDEV�n������̏ޏ ����&�8�J�\�n� ��������ȟڟ���>�PALT�=7� c_�_�q��������� ˯ݯ���%�7�I��[�m������%�GRI�e۱O����� '�9�K�]�oρϓϥ� �����������#�5�G�ɿ��R�=��Y� �߹���������%� 7�I�[�m������������m�PREG ;�$����K�]�o��� �������������� #5GYk}����$ARG_KPD ?	������  �	$�	[��]���� S�BN_CONFIQG� �%!$"�CII_SAVE  �D;� �TCELLSET�UP 
�
%  OME_IO���%MOV_H8���REP�����UTOBACK�s�	AFRwA:\� �,�^'`� �<(�� M+@ �23/04/�01 14:33:48���/0�/�/�/-,��?/?@A?S?e?w?�?��? �?�?�?�?�?O�?5O GOYOkO}O�O�O,O�O �O�O�O__�OC_U_�g_y_�_�_�_�Ё � (!_#_\AT�BCKCTL.T�MP DATE.D:��_oo,o>o#�INI:�o%7~#MESSAGS�]a^� hkODE_AD�V7G�eO����o#PAUS�a!��� ,,		�� ��ow �o-9;M�q ���������;����d�`TSK�  �m</Bo UgPDT�`[gd����fXWZD_ENqB[d3��STAZe�����WEPLS�CH R+   b��.�@� R�d�v���������П �����*�<�N�`� r���������̯ޯ�����RODނ2.�4���/��>� %V�{������� ÿտ�����/�A��SϾWEROBGRP`��r�GWEWEL �2�D� ��h�����'�9�K� ]�o߁ߓߥ߷��߼	�XIS%UN��8�D��� 	r�� ��@�+�d�O��s���������MET�ER 2b�_ �P��&���J���SC�RDCFG 1v�! �[[?�������������5/�
QW��M_ q����2� %7I���!GR�Р��o��PNAME 	��s	$�_EDY`�1s�� 
 ��%-�PEDT- v��/*/j�� �����.��µ���X��/:����%2�/ ���/a/��G(�//?v/�/?�/�#3g?�/�? �/>�?�?B?T?�?x?�#43O�?�O�?>\O@�OO O�ODO�#5�O oOL_�O>(_�_�O�O�__�#6�_;_o__ >�__o�_�_No�_�#7�oo�o+o>�o+ ro�o�o�#8c/�//�=��>P�t�#9/��|���=X�Ï
����@��!CR�/�oG�Y�} "���ԏ�|�
���?NO_DEL���GE_UNUSE���IGALLO�W 1��  � (*SYS�TEM*��	$S�ERV_u�.�G�P�OSREGP�$8r�.�G�NUMu������PMU����LAY��.��PMPALTǧCOYC10Ԟ�Ѡ<ծ�ULSUǯ����r���L#�\�B�OXORIy�CU�R_I���PMC�NVæI�10�����T4DLIB�@�b�	*PROG�RAO�PG_cMIծ���ALߵ����B<�G��$FLUI_RECSU�u��j�������������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r�������������e��LAL_OUT 6��q#�WD_ABO�R��i�ITR_�RTN  �����l�NONSTO���� ��CCG�_CONFIG �7�7���8������E_RIA_�I���, ����FCFG ����5_LImM^�2� � 	n���<�j�ߥ蜀�dP}AV�GP 1?��-�?�C�� C��  C�b�fԪb�f�f�b��f0�D`�DD���
��4���Dv�DZlT~����Vx�D/�9�C��M�W�a��?����HE��u�"G�_P��1�  ��d/v/�/�/�/��/�/HKPAU�Sf�16�,  ���/ ?6�?L?2?\? �?h?�?�?�?�?�?�?�O�?6OHO.OlO
O�9?��h�CO�LLECT_90s	`�N�GEN߰���~��B�ANDE�C�s���12�34567890�!W��a�O_1V��
 H+���)l_�_a� k_}_�_b��_�_o�_ �_	obo-o?oQo�ouo �o�o�o�o�o�o: )�M_q��@�����Fm�K� �N�FIO !
Y�A��������ظ�ʏb�TR� 2"F�(��}�
�؎���#q�� %[�_MkORm$� �) ���������ǟ���Pٛd��n%r�, %I?	!	!�>���KH�*��$R9&�Ow��v�v�C4  A�l�
� x��AA��Cz  B�fPB}���C  @��������:d�U
\�IS'f�\��T_DEF*� ��%�+�����IN�US�&,@�KEY_TBL  ��,v� �	
��� !"#�$%&'()*+�,-./*W:;<=>?@ABC��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~�����������������������������������������������������������������������������������������������������������������������������������������6�d�L�CKI���d�I�ST�As�>�_AUTO�_DO��m���I�ND�D�δAR_T1�Ͽ�T2��������A�XC� 2(�q�cP8
SONY XC-56{��u��U��@����� ��А~�HR5XY ���έ�R57����ACff���6�H� $� m��Z�������� ���!���E�W�2�{�܍��TRL�LE�TE!��T_S�CREEN ~�
kcsc"�UD�MMENU �1)�	  <u��1�:o `CLr����� �� &_6H �l~����/ ��I/ /2//V/h/ �/�/�/�/�/�/�/3? 
??B?{?R?d?�?�? �?�?�?�?�?/OOO eO<ONO�OrO�O�O�O �O�O_�O_O_&_8_ ^_�_n_�_�_�_�_o �_�_oKo"o4o�oXo jo�o�o�o�o�o�o�o�5+���_MANU3ALH��DB9�0������DBG_ER�RL�*����C >���~uq�NUMLIM���dn�ޠDBPXWORK 1+���L�^�p�������DBTB_�� Q,�}����u�RqDB_AWAY}s�͡GCP n�=s����_AL
����yrYGл�n�nx�_�p 1-q�
́.�
;�y�z�g�l����_M��IS�����@A���ONTImM���n��ޖ�4�
X�I�MOTN�ENDM�H�REC�ORD 13��� �����G�O� t�b���������į֯ m�ޯ�t�)���M�_� q������˿:�� ��%���Iϸ�m�ܿ �ϣϵ���6���Z�� ~�3�E�W�i��ύ��� �� ��������z�/� ��:���w����� ��@���d��+�=�O����s�^�l�����Oi������b�M��sN��������[���);�_JX���W�����N/��9/�k0�.:/q/�/���TO�LERENC��B��>��L��upC�SS_CNSTC�Y 24,���p�/<���/??(?>? L?^?p?�?�?�?�?�? �?�? OO$O6OHO�$�DEVICE 25�+ І�O�O �O�O�O�O__+_=_�O_���#HNDGDg 6�+ՀCzi^_LS 27�Ma_ �_�_�_oo'o9oc_��"PARAM �8U�%�duKd�$SLAVE 9�]�nW_CFG :�koKcdMC:�\� L%04d.'CSVJo<�c�ofr6+"A sCHp�QA��Kn*_}g�Kf�Or|q�zyyq�`�JPѬsk~<�ρ��lRC_OUT �;�MρOo_SG�N <K�4����mE15-A�PR-23 11�:32p�a0=13�4:35p�F V�t�g��c�Knd�+�@�S�Þ�j�x��z��cVERSIO�N �V�4.0.1��EF�LOGIC 1=^�+ 	�x�`���q��PROG�_ENB)��V2�U�LS� �V�_�ACCLIM����c�q�WRSTJNɐ�3��a��MO;�uq�b��I?NIT >�*K�v�a ��OPT�`� ?	�Ȓ
 ?	R575Kc��74!�6"�7"�50F�ׄL�2"��xp�|އ��TO  ��z�ů߆V֐DEXҞ�d&��pݣPA�TH A�A�\˯*�<��+HCP�_CLNTID y?�c �{�G#|��!IAG_G�RP 2C�i Q�	��ؿÿ���� ��Dϒ�m�p1m10 89�012345678n���=�� ?Ϝ� �ω������r��� ���!�3���\�n����q�Gߩ߻ߙ��� ��{����9�K�)�o� ���U�g�������� �����3�Y�7�i��� �+�u������� ��/gyW�� 9���	�-? �>χ:ϫ�� ��|���;/&/_/�˰_O 4Q/�/A/ #�/g�/?!?혒$ -?W?�/g?�?o?�?�? m�?E/O�?ODO/O hOSO�OwO�O�O�O�O��O
_�O.__R_��<�p c_�_�_ C_�_�_�_�_�_o0o �_@ofoQo�ouo�o�o��o��CT_CON�FIG D��|ʓ]�eg�u���STBF_TTS��
J�)s��}�xq:<v�pMAU��?�~Q�MSW_CF�`�E��  ��OCoVIEWPpF�}�a�������� *�<����e�w����� ����N������+� =�̏a�s��������� ͟\����'�9�K� ڟo���������ɯX� ����#�5�G�Y�� }�������ſ׿f������1�C�Uϡ|RC�sG]r!�c΍� �ϱ�����
���.�t�SBL_FAUL�T H�ʥxH�G�PMSK2w[��`TDIAG Iy�qUt��UD�1: 6789012345��x��c�P�o����*�<� N�`�r�������@������;�Vp����@8r��\��fTRECP�ߣ�
�ԣ��� ��������1C Ugy��������	0�B�?f�U�MP_OPTIO1N2pT�aTR�r3s:X��PME1uu�Y_TEMP  È�3B�Vp���A��UNI�np4u���YN_B�RK J��bE�DIT_y�ENT� 1K��  �,&MAIN_�SOLDADUR�AOP&	G#O�N L/P&IR?_HOME v/5��&REQMEN�U�/�/�?r� �/-??Q?8?`?�?n? �?�?�?�?�?O�?)O ;O"O_OFO�OjO|O�O �O�O�O�O_�O7__�[_m_T_�_xY MG?DI_STA��ql�%NC�S1L�{� ��_�_P
Pd7Yoko}o�o�o �o�o�o�o�o1 CUgy���� ����� �.�Fa .�T�f�x��������� ҏ�����,�>�P� b�t���������6�� ����#�=�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������۟���	�� 5�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߹�ӿ ������-�#�I�[� m����������� ���!�3�E�W�i�{� �������������� ��7�ASew�� �����+ =Oas����� ����///9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?��?�?�? O'/1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �?�_�_�_oOo;o Mo_oqo�o�o�o�o�o �o�o%7I[ m���_��� �o)o3�E�W�i�{� ������ÏՏ���� �/�A�S�e�w����� ��џ����!�+� =�O�a�s��������� ͯ߯���'�9�K� ]�o��������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ��������� ��1�C�U�g�yߋ� �߷����������� -�?�Q�c�u���� ����������)�;� M�_�q������ߝ��� ����	���%7I[ m������ �!3EWi{ ��������� ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?���? �?�?�?/O'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�?�_�_�_�_O oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��_� ����_��)�;� M�_�q���������ˏ ݏ���%�7�I�[� m�������ǟٟ� ��!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� =�O�a�sυϗϩϻ� ��������'�9�K� ]�o�鿛��߷����� �����#�5�G�Y�k� }������������ ��1�C�U�g�y��� ������������	 -?Qcu��� ����); M_q��y��� ���//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?� ��?�?�?y?��?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_O_a_{?�?�_�_�_ �_�?�_oo'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk �_�����_�� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�}������ ���ɟ���)�;� M�_�q���������˯ ݯ���%�7�I�[� u�g�������ϟ�� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�m���ߛ� �߿�ٿ������+� =�O�a�s����� ��������'�9�K� ��w߁����������� ����#5GYk }������� 1CUo�y� �������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?gU?�?�?�?��? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O��O_!_3_E__? ��$ENETMOD�E 1M�5��  o0�o0j5�_�[nPRR�OR_PROG %{Z%i6�_�Y�U�TABLE  {[�?-o?oQo_g�R�SEV_NUM ��R  ���Q�`�Q_AUTO_ENB  �U܃S�T_NO�a �N{[�Q�b  �*��`��`��`��`�`+�`�o�d�HIS}cm1�P�k_�ALM 1O{[� �j4�li0+ �������_vb�`  {[��a�R2�nPTCP_�VER !{Z!��_�$EXTLO�G_REQ3v蜩i��SIZ���SkTK���e􁂿TOL  m1D�z;r�A �_BWD�瀠f��Rv��DI� P�5���Tm1�S�TEP)�;�nPU�O�P_DȌlQFD�R_GRP 1Q{Y�ad 	-�ʟ�P����E%����?�#���[��� �
� �������� !��D�/�h�S���w� �������ѯ
���.��W
$�]�fvM����x������B�  ��A�  @�338��UO��Ϳ���9�$�F�6 F@]�[�g�"σ�F�? ?�  �Ϙ��<P���;O���9 n���r��������K����/ 舡�[������[�FEATURE �R�5��Q�ArcTool� D�m2Eng�lish DictionaryO��4D Stand�ardH�Anal�og I/OG�A�Z�e Shift���rc EQ P�rogram S�elect��So�ftpar����W�eld��cedu�res��@�Cor�e��?�Rampi�ng��uto��w�a'�Update�M�matic B�ackupM�{�g�round Ed�itE�R�Came�ra��F��Cel�l�ܠ�nrRnd�Im���ommo�n calib 3UI����sh����b�c&�.���neCӖ.�ty��s����n����Monito�rb�ntr>�el�iab��N�DHC�PD۷�ata A�cquis���iagnosw�����ocument �Viewe���u�a#�heck S�afety	�R�h{an� Rob��rv��qF
�N�k�s" F��(�R�xt� weavx�ch�J�xt. DIO�$�nfiG� en]dS Err��L���s�	r���  ��L�FCTN M�enu; �  TPw Infac(�R�Gen��l�E�q L�]��p �Mask Exc�O g�HTJ��x�y Sv#�ig�h-SpeS Sk�i����$�mmu�nicv�on�Hour1����M�conn}�2(n{crLstruc��M�KAREL C�md. L�ua��E#Run-Ti�� Env;(_�+�z�sx�S/WO�L?icense5"�� Book(Sy�stem)L�MA�CROs,�/O�ffse�MMR�����MechStop��t�����%i���6xS ��x�v1>od��wit��T8����.$�r;Op�tm�?�#��fil�"�'g��%ult�i-T�E�P�PC�M fun4'�9o���6E�MRegi�� r��6ri F
KRF��Nu����nH��Adju�hN��<�٦MtatuNA�O�
Q�RDMUot>`�scovei��Eem0�nw��ER8Z� ^ues��9W�o$�_0N�SNPX� b�"H�SNJCCli}^��urh�D�_z� %4ujUo� =t1ssagE�jU�A�{_F� U��!n�/IKeMILI�B;obP Fir�m^�%nP1Acc<����TPTX��deln� XoaA��%�&morIP SimGula����fu� AP]�j���3&��gev.eV�ri3 ��oUSB po,���iP� a bunexceptS `P(Dbu�uVC�r��8V���rvoh�u�[�{S�PSC�e.
�SUIK�W� �8<�b Pl�FX�Z ���M�#��FQ�uvn�ԇGri=d
Qplay΍"`���R�r.wڊ�R�C�g�100iD�/1450��la�rm Cause�/Pedj�Asc{ii��Load" �v�Upl����yc���k"Y@Pp@ %RA�p��l�"�NRTL��oS�Online Hel���6L�6�L@IA�trG�64MB DRAM��N\�FROe���tl!:�0.L�mai#��[:�L%�Supmr�1pNIР� �cro�L`S�U��V�Rmi܉F�vrt2SK���� ��W�i�������̿ÿ տ����%�/�\�S� eϒωϛ��Ͽ����� ���!�+�X�O�aߎ� �ߗ��߻�������� �'�T�K�]���� ������������#� P�G�Y���}������� ��������LC U�y����� ��H?Q~ u������� //D/;/M/z/q/�/ �/�/�/�/�/�/	?? @?7?I?v?m??�?�? �?�?�?�?OO<O3O EOrOiO{O�O�O�O�O �O�O__8_/_A_n_ e_w_�_�_�_�_�_�_ �_o4o+o=ojoaoso �o�o�o�o�o�o�o 0'9f]o�� ������,�#� 5�b�Y�k�������Ώ ŏ׏���(��1�^� U�g�������ʟ��ӟ ���$��-�Z�Q�c� ������Ư��ϯ��  ��)�V�M�_����� ��¿��˿���� %�R�I�[ψ�ϑϾ� ����������!�N� E�W߄�{ߍߺ߱��� �������J�A�S� ��w��������� ���F�=�O�|�s� ������������ B9Kxo�� �����> 5Gtk}��� ��/�/:/1/C/ p/g/y/�/�/�/�/�/  ?�/	?6?-???l?c? u?�?�?�?�?�?�?�? O2O)O;OhO_OqO�O �O�O�O�O�O�O_._ %_7_d_[_m_�_�_�_ �_�_�_�_�_*o!o3o `oWoio�o�o�o�o�o �o�o�o&/\S e������� �"��+�X�O�a��� ���������ߏ�� �'�T�K�]������� �����۟���#� P�G�Y���}������� �ׯ����L�C� U���y�������ܿӿ ��	��H�?�Q�~� uχϡϫ�������� ��D�;�M�z�q߃� �ߧ�������
��� @�7�I�v�m���� ����������<�3� E�r�i�{��������� ����8/An ew������ �4+=jas �������/ 0/'/9/f/]/o/�/�/ �/�/�/�/�/�/,?#? 5?b?Y?k?�?�?�?�? �?�?�?�?(OO1O^O UOgO�O�O�O�O�O�O��O�O$_Q  ?H541S?Q�2DVR782EW5�0EUJ614iW7�6EUAWSPQW1��WRCRuX8�VT=U�VJ545iX�V�VCAMEUCLI�O�VRI�WUIFzQV6�WCMSCh^�VSTYLiW2�VoCNREQV52�VwR63PWSCHEU�DOCVqfCSU�EUORS�VR86�9iW0tW88DVE�IOfR54\VR{69�VESET�W��WJ�YWMGEUM�ASKEUPRXY�5h7EVOC�V�`3`�X\V�`hXgX53�f�H^xLCHvOP�LvJ50HvPSƛwMC�W�p�g55�tVMDSW�w;wOP;wMPR�Va`0v\�`hVPCMg0�l�`tW50�51�W�51P�0�VPRSv�g690vFRD�V�RMCN)f�hH9=3hVSNBAg_w/SHLB)fM߇a`�XgNNlx2hVHTC�VTMI4fYP�f�TPAfTPTXF�EL���p�g8[W�YPDVJ95�VTU�T<w950vUEC�vUFR�VVCC���O�VVIP4fC�SCL��`I�xtVW�EB�VHTT�W6nWgWIO��CG�{IG�IPGS=��RC4fHZXR66V�VR7�gRN�2HvRjz40vu�tV`DV�NVD�fD0��Fn�CTO�WNN0v�OL'hENDQVL�×SLM�fFVR e XK�]�o������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U� g�yߋߝ߯������� ��	��-�?�Q�c�u� ������������ �)�;�M�_�q����� ����������% 7I[m��� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-?Qcu �������� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�e� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ����������'�  H�541)�C�2H�R�782I�50I�J�614y�76I�A�WSPY�1��RC�R��8��TU��J�545yܘ�VCA�MI�CLIO�R]I�UIFY�6���CMSCY��ST�YLy�2��CNR�EY�52��R63�X�SCHI�DOC�V��CSUI�OR�S��R869y�0v��88H�EIOh�wR54h�R69��OESET�۷�J���WMGI�MASK^I�PRXY��7I�OC(��3��hڅ�x�w�53�HL�CH��OPL��J�50��PSgMCا�u ��55��MD�SW���OP��M�PR(�����%�x�P�CMH�0����5m051��51X�0��PRSx�69���FRD�RMC�Ny��H93x�S�NBAI�SHL�By�M+���NN�(2x�HTC��T�MI��e��TPA�h�TPTXi*EL��u �8g�e�H�J�95��TUT��9�5��UEC��UF]R�VCC8<O��wVIP��CSC�*r��Ii��WEB���HTT��6��WImO�:CG�;IG�;oIPGS�:RC���Hf�R66��R7�g�RV2��R&4���5@��U�H�NVD�x�D0�KF�LCTmO��NN��OLw��ENDY�LG;SLMx�FVRh�(�O_ a_s_�_�_�_�_�_�_ �_oo'o9oKo]ooo �o�o�o�o�o�o�o�o #5GYk}� �������� 1�C�U�g�y������� ��ӏ���	��-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭߿� ��������+�=�O� a�s��������� ����'�9�K�]�o� ���������������� #5GYk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ����������%�1�S�TD,�LANGM�H�`�r߄ߖߨ� ����������&�8� J�\�n������� �������"�4�F�X� j�|������������� ��0BTfx ������� ,>Pbt�� �����//(/�:/L/^$RBTL�OPTNu/�/�/�/�/�+DPNK��/�/? ?/?M�$�S?e?w?�? �?�?�?�?�?�?OO +O=OOOaOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�_�_�_�_�_ �_�_�_o#o5oGoYo ko}o�o�o�o�o�o�o �o1CUgy �������	� �-�?�Q�c�u����� ����Ϗ����)� ;�M�_�q��������� ˟ݟ���%�7�I� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O�__99'U��$FEAT_AD�D ?	����TQ\P  	$Xe_w_�_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o ���������#5GGTDEM�O RTY   $X���� ����///&/8/ R/\/�/�/�/�/�/�/ �/�/�/+?"?4?N?X? �?|?�?�?�?�?�?�? �?'OO0OJOTO�OxO �O�O�O�O�O�O�O#_ _,_F_P_}_t_�_�_ �_�_�_�_�_oo(o BoLoyopo�o�o�o�o �o�o�o$>H ul~����� ��� �:�D�q�h� z�������ݏԏ�� 
��6�@�m�d�v��� ����ٟП���� 2�<�i�`�r������� կ̯ޯ���.�8� e�\�n�������ѿȿ ڿ����*�4�a�X� jϗώϠ�������� ���&�0�]�T�fߓ� �ߜ������������ "�,�Y�P�b���� �����������(� U�L�^����������� ������ $QH Z�~����� �� MDV� z������� //I/@/R//v/�/ �/�/�/�/�/�/?? E?<?N?{?r?�?�?�? �?�?�?�?
OOAO8O JOwOnO�O�O�O�O�O �O�O__=_4_F_s_ j_|_�_�_�_�_�_�_ oo9o0oBooofoxo �o�o�o�o�o�o�o 5,>kbt�� ������1�(� :�g�^�p�������ӏ ʏ܏�� �-�$�6�c� Z�l�������ϟƟ؟ ���)� �2�_�V�h� ������˯¯ԯ��� %��.�[�R�d����� ��ǿ��п���!�� *�W�N�`ύτϖ��� ����������&�S� J�\߉߀ߒ߿߶��� ������"�O�F�X� ��|���������� ���K�B�T���x� ������������ G>P}t�� ����C :Lyp���� ��	/ //?/6/H/ u/l/~/�/�/�/�/�/ ?�/?;?2?D?q?h? z?�?�?�?�?�?O�? 
O7O.O@OmOdOvO�O �O�O�O�O�O�O_3_ *_<_i_`_r_�_�_�_ �_�_�_�_o/o&o8o eo\ono�o�o�o�o�o �o�o�o+"4aX j������� �'��0�]�T�f��� ������������#� �,�Y�P�b������� ����������(� U�L�^����������� �ܯ���$�Q�H� Z���~��������ؿ ��� �M�D�Vσ� zόϦϰ�������� 
��I�@�R��v߈� �߬���������� E�<�N�{�r���� ���������A�8� J�w�n����������� ����=4Fs j|����� �90Bofx �������/ 5/,/>/k/b/t/�/�/ �/�/�/�/�/?1?(? :?g?^?p?�?�?�?�? �?�?�? O-O$O6OcO ZOlO�O�O�O�O�O�O �O�O)_ _2___V_h_ �_�_�_�_�_�_�_�_ %oo.o[oRodo~o�o �o�o�o�o�o�o! *WN`z��� ������&�S� J�\�v���������� ڏ���"�O�F�r�  i����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(:�L^p   qk������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ���������&� 8�J�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x��������������� ,>Pbt� ������ (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�_�_�_oo&o 8oJo\ono�o�o�o�o �o�o�o�o"4F Xj|����� ����0�B�T�f� x���������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*�<�N�`�r��� �����������&� 8�J�\�n��������� ��������"4F Xj|����� ��0BTf
vzm��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n���� �����������"�4� F�X�j�|��������� ������0BT fx������ �,>Pbt �������/ /(/:/L/^/p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\n��� ������"�4� F�X�j�|�������ď ֏�����0�B�T��f�x��$FEAT�_DEMOIN [ {�����~�}��INDEX��������ILEC�OMP S�;��ޑ�����ԐSETUP2 �Tޕ���  N �ѓ_A�P2BCK 1U~ޙ  �)y�DG�V�%=�z�~�� h���{�<�ѯ`����� �+���O�ޯs���� ��8�Ϳ߿n�ϒ�'� 9�ȿ]�쿁�ώϷ� F���j���ߠ�5��� Y�k��Ϗ�߳���T� ��x����C���g� �ߋ��,���P����� �����?�Q���u�� ��(�����^����� )��M��q�� 6��l�%� 2[���D �h�/�3/�W/ i/��//�/@/�/�/ v/?�//?A?�/e?�/ �?�?*?�?N?�?�?�? O�?=O�?JOsO�!��P%� 2:�*�.VRzO�O2@*��O�O/C�O_E�@P�C_H_2@FR6�:3_t^_�_'[T ���_�_]U�_�\���_<o F*.F�OOo"1A	_S=o|lo�o/kSTM�o�o\RbPD�o }�o$/kH�o�W�gE�0jGIF���e���-�0jJPG7�a��e`M�
����(ZJS����2@w�ҏ��%
�JavaScri3pt�;�CS�h���fU�� %Ca�scading �Style Sh�eets��@
A�RGNAME.D)Tß&L�`\ן�������ğ�DISP*���`[����*�����H�
TPEINS.XML˯�w�:\߯����Cu�stom Too�lbar �O�PA?SSWORD��$N?FRS:\c�"�� %Passw�ord Config���?�|��#� YOG�ֿk�}�ϡ�0� ����f��ϊ�߮��� U���y��r߯�>��� b���	��-��Q�c� �߇���:�L���p� �����;���_���� ��$���H�����~� ��7����m���  ��V�z!� E�i{
�.� Rd��/�/S/ �w//�/�/</�/`/ �/?�/+?�/O?�/�/ �??�?8?�?�?n?O �?'O9O�?]O�?�O�O "O�OFO�OjO|O_�O 5_�O._k_�O�__�_ �_T_�_x_oo�_Co �_go�_o�o,o�oPo �o�o�o�o?Q�o u��:�^� ��)��M��F��� ���6�ˏݏl���� %�7�Ə[���� � ��D�ٟh�ҟ���3� W�i��������ï R��v������A�Я e���^���*���N�� ����Ϩ�=�O�޿s� ϗ�&�8���\��π� ��'߶�K���o߁�� ��4�����j��ߎ�#�����Y�;��$FI�LE_DGBCK� 1U��F���� <� �)
SUMM?ARY.DGc��OMD:������Diag Su�mmary����
CONSLOG�������[���Co�nsole lo�g\���	TPACCNQ���%�������TP Acco�untin}����FR6:IPKD?MP.ZIP��
'`����Exc?eptiond���MEMCHEC�K��8����o�M�emory Da�ta�;�/YF)	FTPN�?��C�q�mmen�t TBDl;�L� =�)ETHERNETa������Ethe�rnet s�fi�gura���VDCSVRF`FX�q/�%6  v�erify alylt/>�M+�1%DIFFi/O/a/�/�� %�(dif�f�/�'�6 CHG01�/�/�/{?�!?,�?�"*f992q?X?@j?�?
?�?�?@23�?8�?�?�O O�O�9FVTRNDIAG.LS�O`OrO�_��A ��no�stic_>�T6�a)UPDA�TES.MP3_��FRS:\K_�]���Updates� List�_�P�SRBWLD.C	M�_�wR�_�_p��PS_ROBOW�EL����AHADOW�O�O�O�o��Shadow Changes�o�qQbNOT�I;/lo~o�N?otific"�o;�+@AG��j� �9�����w� ��B��f�x���� +���ҏa�������� '�P�ߏt������9� Ο]�����(���L� ^�ퟂ����5���ܯ k� ���$�6�ůZ�� ~������C�ؿ�y� ϝ�2���?�h����� ϰ���Q���u�
�� ��@���d�v�ߚ�)� ��M����߃���<� N���r����7��� [������&���J��� W������3�����i� ����"4��X��| ��A�e� �0�Tf�� ��O�s//� >/�b/�o/�/'/�/ K/�/�/�/?�/:?L? �/p?�/�?�?5?�?Y? �?}?�?$O�?HO�?lO ~OO�O1O�O�OgO�O �O _2_�OV_�Oz_	_ �_�_?_�_c_�_
o�_ .o�_Rodo�_�oo�o �oMo�oqo�o< �o`�o��%�I ����8�J�� n����!���ȏW�� {��"���F�Տj�|� ���/�ğ֟e����� ���+�T��x���� ��=�үa������,� ��P�b�񯆿���9� ���o�ϓ�(�:�ɿ ^��ϔ�#ϸ�G��� ��}�ߡ�6���C�l��N��$FILE_�FRSPRT  ���V�������MDO?NLY 1U��N�� 
 �)�MD:_VDAEXTP.ZZZs��$���
�6%�NO Back �file ��N�S�6�\��߀�I� �������i������ 4���X�j������� ��S���w���B ��f����+�O ����>P� t�'��]� �/(/�L/�p/�/�/�/5/�/�/��VI�SBCK�؝����*.VD�/'?� �FR:\� ION?\DATA\?�"�� Vision VD(�S?a/�? �?�/�?�/�?�?O+O �?OO�?sO�OO�O8O �O\OnO_�O'_9_�O ]_�O�__�_�_F_�_ j_�_o�_5o�_Yo�_ �_�oo�o�o�o�oxo �oC�og�o� �,�P�t���{�LUI_CON�FIG V���	1&� $ ���{��}�������0ŏ׏�e�|x�� !�3�E�W�g������� ����ҟi����,� >�P��t��������� ίe����(�:�L� �p���������ʿa� � ��$�6�H�߿l� ~ϐϢϴ���]����� � �2�D���h�zߌ� �߰���Y�����
�� .���?�d�v���� C���������*��� N�`�r�������?��� ����&��J\ n���;��� �"�FXj| ��7����/ /�B/T/f/x/�/!/ �/�/�/�/�/?�/,? >?P?b?t?�??�?�? �?�?�?O�?(O:OLO ^OpO�OO�O�O�O�O �O _�O$_6_H_Z_l_ ~__�_�_�_�_�_�_ �_ o2oDoVohozoo �o�o�o�o�o}o�o .@Rd�o��� ���y��*�<� N�`����������̏ ޏu���&�8�J�\� 󏀟������ȟڟq� ���"�4�F�X��|�@������į֯f���|�$FLUI_�DATA W������j���RESUL�T 2X�0�� �T�/w�izard/gu�ided/ste�ps/Expert�g�y����������ӿ���	��)���Continue with GD�ance)�d�vψ� �ϬϾ���������*� �-��I�0 �r�I�	�l�i��;�ps,� ����������� �2� D�V�h�z�9�r���� ����������1�C� U�g�y���i�[�m��}��torch�� %7I[m �������� !3EWi{�� ������������wproc��U/g/ y/�/�/�/�/�/�/�/ 	??�??Q?c?u?�? �?�?�?�?�?�?OO@)O��DO/�����M�TimeUS/DST3O�O�O�O�O __'_9_K_]_o_2�DisablR� �_�_�_�_�_�_o"o�4oFoXojo|n�j�eOWOiO{O�O�B24�O/AS ew����~_�_ ���+�=�O�a�s� ��������͏�o�o�o��o��:�L�RegionЏ_�q����������˟ݟ���.�AmericaI/ M�_�q���������˯@ݯ���.�ہyE����]��1��BEdi ��$���ſ׿������1�C�U�g�*; T�ouch Pan�el �� (re�commen��) uϺ���������&� 8�J�\�n�-��=�O���s����Bacces<���*�<�N�`��r�����)<C�onnect t�o Network�� ��$�6�H�Z��l�~���������1��0鏣����!�ߝ@�IntroductK�^p���� ��� -?6H Zl~�����0��/ / =O�� =/�b0�/�/�/�/ �/�/�/?#?5?G?Y? k?*�?�?�?�?�?�? �?OO1OCOUOgO׈�@ ]/G*���~�O�O}/�O�O__ *_<_N_`_r_�_�_�_ �_y?�_�_oo&o8o Jo\ono�o�o�o�ouO �O�O�O�O4FX j|������ ���_0�B�T�f�x� ��������ҏ���� ��o�o�o_�!���� ����Ο�����(� :�L�^���������� ʯܯ� ��$�6�H� Z�l�+�=�O���s�ؿ ���� �2�D�V�h� zόϞϰ�o������� 
��.�@�R�d�v߈� �߬߾�}��ߡ��ſ *�<�N�`�r���� ����������%�8� J�\�n����������� ��������1��U �|������ �0BTf%� �������/ /,/>/P/b/!�/E �/ik/�/�/??(? :?L?^?p?�?�?�?�? w�?�? OO$O6OHO ZOlO~O�O�O�Os/�O �/�O_�?2_D_V_h_ z_�_�_�_�_�_�_�_ 
o�?.o@oRodovo�o �o�o�o�o�o�o�O _�O3]_��� ������&�8� J�\�o��������ȏ ڏ����"�4�F�X� a;����q֟� ����0�B�T�f�x� ������m�ү���� �,�>�P�b�t����� ��i�{������ß(� :�L�^�pςϔϦϸ� ������ ߿�$�6�H� Z�l�~ߐߢߴ����� �����Ϳ߿�S�� z������������ 
��.�@�R��v��� ������������ *<N`�1�C� g����&8 J\n���c�� ���/"/4/F/X/ j/|/�/�/�/q�/� �/�?0?B?T?f?x? �?�?�?�?�?�?�?O ?,O>OPObOtO�O�O �O�O�O�O�O_�/%_ �/I_?p_�_�_�_�_ �_�_�_ oo$o6oHo ZoO~o�o�o�o�o�o �o�o 2DV_ w9_�]__��� 
��.�@�R�d�v��� ����koЏ���� *�<�N�`�r������� gɟ����Ï&�8� J�\�n���������ȯ گ�����"�4�F�X� j�|�������Ŀֿ� �����ݟ'�Q��x� �ϜϮ���������� �,�>�P��t߆ߘ� �߼���������(� :�L��U�/�y��e� ������ ��$�6�H� Z�l�~�����a����� ���� 2DVh z��]�o���� ��.@Rdv� ��������/ */</N/`/r/�/�/�/ �/�/�/�/?��� G?	n?�?�?�?�?�? �?�?�?O"O4OFO/ jO|O�O�O�O�O�O�O �O__0_B_T_?%? 7?�_[?�_�_�_�_o o,o>oPoboto�o�o WO�o�o�o�o( :L^p���e_ ��_��_�$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� ���=��d�v��� ������Я����� *�<�N��r������� ��̿޿���&�8� J�	�k�-���Q�S��� �������"�4�F�X� j�|ߎߠ�_������� ����0�B�T�f�x� ���[Ͻ������� �,�>�P�b�t����� ������������( :L^p���� ���������E �l~����� ��/ /2/D/h/ z/�/�/�/�/�/�/�/ 
??.?@?�I#m? �?Y�?�?�?�?OO *O<ONO`OrO�O�OU/ �O�O�O�O__&_8_ J_\_n_�_�_Q?c?u? �?�_�?o"o4oFoXo jo|o�o�o�o�o�o�o �O0BTfx ��������_ �_�_;��_b�t����� ����Ώ�����(� :��o^�p��������� ʟܟ� ��$�6�H� ��+���O���Ưد ���� �2�D�V�h� z���K���¿Կ��� 
��.�@�R�d�vψ� ��Y���}��ϡ��� *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n������� ��������1���X� j�|������������� ��0B�fx ������� ,>��_!��E� G����//(/ :/L/^/p/�/�/S�/ �/�/�/ ??$?6?H? Z?l?~?�?O�?s�? �?�/O O2ODOVOhO zO�O�O�O�O�O�O�/ 
__._@_R_d_v_�_ �_�_�_�_�_�?�?�? o9o�?`oro�o�o�o �o�o�o�o&8 �O\n����� ����"�4��_=o oa���Mo��ď֏� ����0�B�T�f�x� ��I����ҟ���� �,�>�P�b�t���E� W�i�{�ݯ����(� :�L�^�p��������� ʿܿ�� ��$�6�H� Z�l�~ϐϢϴ����� �ϩ���ͯ/��V�h� zߌߞ߰��������� 
��.��R�d�v�� ������������ *�<����߁�Cߨ� ��������&8 J\n�?��� ���"4FX j|�M��q���� �//0/B/T/f/x/ �/�/�/�/�/�/�? ?,?>?P?b?t?�?�? �?�?�?�?�O�%O �LO^OpO�O�O�O�O �O�O�O __$_6_�/ Z_l_~_�_�_�_�_�_ �_�_o o2o�?SoO wo9O;o�o�o�o�o�o 
.@Rdv� G_������� *�<�N�`�r���Co�� goɏۏ���&�8� J�\�n���������ȟ ڟ����"�4�F�X� j�|�������į֯�� ߏ���-��T�f�x� ��������ҿ���� �,��P�b�tφϘ� �ϼ���������(� �1��U��A��߸� ������ ��$�6�H� Z�l�~�=Ϣ������ ����� �2�D�V�h� z�9�K�]�o������� 
.@Rdv� ������� *<N`r��� ���������#/�� J/\/n/�/�/�/�/�/ �/�/�/?"?�F?X? j?|?�?�?�?�?�?�? �?OO0O�//uO 7/�O�O�O�O�O�O_ _,_>_P_b_t_3?�_ �_�_�_�_�_oo(o :oLo^opo�oAO�oeO �o�O�o $6H Zl~����� �o�� �2�D�V�h� z�������ԏ�o�� �o��o@�R�d�v��� ������П����� *��N�`�r������� ��̯ޯ���&�� G�	�k�-�/�����ȿ ڿ����"�4�F�X� j�|�;��ϲ������� ����0�B�T�f�x� 7���[����ߓ���� �,�>�P�b�t��� ����������(� :�L�^�p��������� �����߭���!��H Zl~����� �� ��DVh z������� 
//��%��I/s/5 �/�/�/�/�/�/?? *?<?N?`?r?1�?�? �?�?�?�?OO&O8O JO\OnO-/?/Q/c/�O �/�O�O_"_4_F_X_ j_|_�_�_�_�_�?�_ �_oo0oBoTofoxo �o�o�o�o�o�O�O�O �O>Pbt�� ��������_ :�L�^�p��������� ʏ܏� ��$��o�o i�+������Ɵ؟ ���� �2�D�V�h� '�y�����¯ԯ��� 
��.�@�R�d�v�5� ��Y���}������ *�<�N�`�rτϖϨ� ����ݿ����&�8� J�\�n߀ߒߤ߶��� ���߫��Ͽ4�F�X� j�|���������� ������B�T�f�x� �������������� ��;��_!�#� �����( :L^p/���� ��� //$/6/H/ Z/l/+�/O�/�/� �/�/? ?2?D?V?h? z?�?�?�?�?��?�? 
OO.O@OROdOvO�O �O�O�O}/�/�/�O_ �/<_N_`_r_�_�_�_ �_�_�_�_oo�?8o Jo\ono�o�o�o�o�o �o�o�o�O_�O= g)_������ ���0�B�T�f�%o ��������ҏ���� �,�>�P�b�!3E W��{�����(� :�L�^�p��������� w�ܯ� ��$�6�H� Z�l�~�������ƿ�� �����͟2�D�V�h� zόϞϰ��������� 
�ɯ.�@�R�d�v߈� �߬߾��������� ׿���]�τ��� ����������&�8� J�\��m��������� ������"4FX j)�M�q��� �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/{�/�?�(? :?L?^?p?�?�?�?�? �?�?�? OO�6OHO ZOlO~O�O�O�O�O�O �O�O_�//_�/S_? _�_�_�_�_�_�_�_ 
oo.o@oRodo#O�o �o�o�o�o�o�o *<N`_�C_� �{o����&�8� J�\�n���������uo ڏ����"�4�F�X� j�|�������q�� ߟ	��0�B�T�f�x� ��������ү���� Ǐ,�>�P�b�t����� ����ο���ß� �1�[���ϔϦϸ� ������ ��$�6�H� Z��~ߐߢߴ����� ����� �2�D�V�� '�9�Kϭ�o������� 
��.�@�R�d�v��� ����k������� *<N`r��� �y������&8 J\n����� �����"/4/F/X/ j/|/�/�/�/�/�/�/ �/?���Q?x? �?�?�?�?�?�?�?O O,O>OPO/aO�O�O �O�O�O�O�O__(_ :_L_^_?_A?�_e? �_�_�_ oo$o6oHo Zolo~o�o�o�o�_�o �o�o 2DVh z���o_��_� �_�.�@�R�d�v��� ������Џ����o *�<�N�`�r������� ��̟ޟ���#�� G�	����������ȯ گ����"�4�F�X� �|�������Ŀֿ� ����0�B�T��u� 7��ϫ�o�������� �,�>�P�b�t߆ߘ� ��i���������(� :�L�^�p����e� �ω������$�6�H� Z�l�~����������� ������ 2DVh z������� �����%O�v� ������// */</N/r/�/�/�/ �/�/�/�/??&?8? J?	-?�?c�? �?�?�?O"O4OFOXO jO|O�O�O_/�O�O�O �O__0_B_T_f_x_ �_�_�_m??�?�_�? o,o>oPoboto�o�o �o�o�o�o�o�O( :L^p���� ��� ��_�_�_E� ol�~�������Ə؏ ���� �2�D�U� z�������ԟ��� 
��.�@�R��s�5� ��Y���Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ�c��� ���ϫ��"�4�F�X� j�|ߎߠ߲������� �߹��0�B�T�f�x� ������������� ���;�����t����� ����������( :L�p���� ��� $6H �i+���c�� ��/ /2/D/V/h/ z/�/�/]�/�/�/�/ 
??.?@?R?d?v?�? �?Y�}�?�?�O *O<ONO`OrO�O�O�O �O�O�O�O�/_&_8_ J_\_n_�_�_�_�_�_ �_�_�?�?�?oCoO jo|o�o�o�o�o�o�o �o0B_fx �������� �,�>��_o!o3o�� Wo��Ώ�����(� :�L�^�p�����S�� ʟܟ� ��$�6�H� Z�l�~�����a�s��� 篩�� �2�D�V�h� z�������¿Կ濥� 
��.�@�R�d�vψ� �ϬϾ������ϳ�ů ׯ9���`�r߄ߖߨ� ����������&�8� ��I�n������� �������"�4�F�� g�)ߋ�M߲������� ��0BTfx �������� ,>Pbt�� W��{����//(/ :/L/^/p/�/�/�/�/ �/�/�/�?$?6?H? Z?l?~?�?�?�?�?�? �?�O�/O��?hO zO�O�O�O�O�O�O�O 
__._@_�/d_v_�_ �_�_�_�_�_�_oo *o<o�?]oO�o�oW_ �o�o�o�o&8 J\n��Q_�� ����"�4�F�X� j�|���Mo�oqo��� �o��0�B�T�f�x� ��������ҟ䟣� �,�>�P�b�t����� ����ί௟��Ï� 7���^�p��������� ʿܿ� ��$�6��� Z�l�~ϐϢϴ����� ����� �2���� '���K����������� 
��.�@�R�d�v�� GϬ���������� *�<�N�`�r�����U� g�y�����&8 J\n����� ����"4FX j|������ ������-/��T/f/x/ �/�/�/�/�/�/�/? ?,?�=?b?t?�?�? �?�?�?�?�?OO(O :O�[O/OA/�O�O �O�O�O __$_6_H_ Z_l_~_�_�O�_�_�_ �_�_o o2oDoVoho zo�oKO�ooO�o�O�o 
.@Rdv� ������_�� *�<�N�`�r������� ��̏ޏ�o���o#��o �\�n���������ȟ ڟ����"�4��X� j�|�������į֯� ����0��Q��u� ��K�����ҿ���� �,�>�P�b�tφ�E� �ϼ���������(� :�L�^�p߂�A���e� ���ߛ� ��$�6�H� Z�l�~�������� ����� �2�D�V�h� z��������������� ��+��Rdv� ������ *��N`r��� ����//&/�� ��	}/?�/�/�/ �/�/�/?"?4?F?X? j?|?;�?�?�?�?�? �?OO0OBOTOfOxO �OI/[/m/�O�/�O_ _,_>_P_b_t_�_�_ �_�_�_�?�_oo(o :oLo^opo�o�o�o�o �o�o�O�O�O!�OH Zl~����� ��� ��_1�V�h� z�������ԏ��� 
��.��oO�s�5 ������П����� *�<�N�`�r������� ��̯ޯ���&�8� J�\�n���?���c�ſ ������"�4�F�X� j�|ώϠϲ����ϕ� ����0�B�T�f�x� �ߜ߮����ߑ��ߵ� �ٿ��P�b�t��� �����������(� ��L�^�p��������� ������ $��E �i{?����� �� 2DVh z9������� 
//./@/R/d/v/5 Y�/�/��/?? *?<?N?`?r?�?�?�? �?�?��?OO&O8O JO\OnO�O�O�O�O�O��/�/�/�O_%Q�$�FMR2_GRP� 1Y%U�� �C4 w B��0	 �0�c_u\`PF�6 F@�S�Q�T�J`Sx�_�]`P?�  �_��_<P�a;O?��9 n�e�]�A`+o=kBH]SB�YPX`;a@�33�ce�\�_�o�Y@UO߯a�o�_�o�o�o �o4XC|g����}9R_CF�G ZF[T ���(�:��{NO� FZ
F0�p� u��|RM_C�HKTYP  �6Q�0NPPPP8QRO=M��_MIN���3W�����|`X9P�SSB�s[%U aV��5��
���uTP_D�EF_OW  ��4NS1�IRCO�M��B��$GENOVRD_DO����1o�THR�� �d��du�_ENB�a� u�RAVC�?S\Ӈހ �@�U"���1��?��P�sj �ՑOU*BPbF\x�sXF�nsU<�� �]�ǯq������3C�
YP�YP�%��d��1A@M�?�U�vY��\#�֐SMT?Sc��RP��4��$HOS�TC�r1dFY߀s��?_P MC�4�L�
��6 _ 27.0Z�1C�  e:χϙϫ� ����u��� ��$�G������	anonymousK�yߋߝ�D���� 	�^P���� 8�:�'�n�K�]�o�� ���Ϸ��������� X�5�G�Y�k�}���� �������0���1 CU��y���� ���,�	-?Q ����������� �//)/pM/_/q/ �/�/���/�/�/? ?%?l~�m?�/�? ��?�?�?�?2/O!O 3OEOWOz?�?�/�O�O �O�O�O.?@?R?d?fO S_�?w_�_�_�_�_O �_�_oo+oN_�O�O so�o�o�o�o__&_ :o'n_K]o� Ho>����� Xo5�G�Y�k�}��o�o �o�o�Ώ0��1� C�U��y��������� ��,�	��-�?�Q�����ENT 1e��� P!ڟ��  ����ï��� ���ί/��;��d� ��L���p�ѿ������ �ܿ�O��s�6ϗ� Zϻ�~ϐ��ϴ���� 9���]� �Vߓ߂߷� z��ߞ��������4� Y��}�@��d���� �������C��g��*�QUICC0 t�P�b�����1��������2��c�!ROUTER�d@R�!PC�JOG��!�192.168.�0.10����CA�MPRT�!b�1� +RT}�/A�h�NAME� !u�!RO�BO�S_CF�G 1du� ��Auto�-started^��FTP��;! ͏ϟf/��/�/�/�/ �/o��/??,?O/=? �/t?�?�?�?�?��/ &/8/OL?n/,O]OoO �O�OZ?�O�O�O�O�O "O�O5_G_Y_k_}_�_ ������ʏ_�_BOo 1oCoUogo._�o�o�o �o�o�_xo	-? Qc�_�_�_��o� o���)��oM�_� q������:���ݏ� ��%�l~���� �����ǟٟ���ď !�3�E�W�i������ ��ïկ���@�R�d� A�x�e����������� ��|�����+�N�O� �sυϗϩϻ��� &�8�:��n�K�]�o� �ߓ�ZϷ��������� "ߤ�5�G�Y�k�}�� �����Ϩ����B�� 1�C�U�g�.������ ������x�	-?�Q��_ERR �f�aqPDU�SIZ  ��^����>�WR�D ?%��� � guest����)�;�SCD_GR�OUP 3g, u!�� ��LOA��RE�S�TM� $v�T_�ENBs �TTP_AUTH� 1h� <!�iPendan�GR.���A!KAREL:*R/[/m-KC�/�/�/�z VISION SETk?�/F!??1?w#U?C?m? g?�?�?�?�?�?�>!$CTRL i��;H��
��F�FF9E3�?���FRS:DEFA�ULT`LFA�NUC Web ?Server`JNB !$��	L�O�O�O_�_,_oWR_CONFIG jp��`OqI�DL_CPU_P5C@��B����Pw BH�UMIN�\�x�UGNR_IO�z�����PNPT_SIM_DO�V��[STAL_S7CRN�V �6F�Q�TPMODNTOqLg�[�ARTY�X@�Q�V� %  gx��SOLNK 1k�}�o�o�o�o�o� �bMASTE��Pzi�UOSLA�VE l�AuRAMCACHE0�(bO'!O_CFGr�c�sUO0��r�CYCLq�uy@_?ASG 1maW�
 �)�;�M� _�q���������ˏݏp��{�rNUM�5�	
�rIPo�wRTRY_CN@��R�
�ra_UPD��a�� �r�p�r�nP~u��u�PS�DT_ISOLC�  P{v"�J_23_DSrd.N��OGg1oP{�<��d<�P� #?��R��?�����Q��̯ޯ𯯯�&�8�J�������*�ЮP�qi��PhpEC�so�UKANJI_�*pK�_³� MONG pp;_��y� (�:�L�^�pϒ~"���qa\EF�ŭ���C�L_L�P'�J�İEYLOGGIN�p�u�F���$�LANGUAGE� �FabyD l<�qLG�qr�y^�a ���xu ��e����P���'U0�����;��cM�CH ;��
��(?UT1:\���� ���������!�@3�E�\�i�{��(����lLN_DISP sP�ئ���f��OC4b�RDz�S��A@�OGBOO/K tM�d��>A���k�X�܏��� ������<O�Y���	>F	Q������N�`��O�_BUFoF 1u�me2kE�j�FB�iG� �G>P} t������/�//C/��~DCS� w�{�=���G��/�/�/|�/Z$IO 1x�{G ğ3D��? *?<?N?b?r?�?�?�? �?�?�?�?OO&O:O JO\OnO�O�O�O�O�OZ�%E�PTM�dh� #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo1o�CoUogoyo�o-��BS�EV�����FTYP�_�o�m���RSh���|��F�L 2y=��� �/�������F(TP����b'�NGNAM�6%.�nV$UPS��GIh������f�_LOA�DPROG %���%	T_ARC�WEL�����MA?XUALRM'��A85�̀l�_PRh���� E�	ˀC��z�M�������,�P �2{� ت	Z�aڀ	�|�f4� �~����������(Ο ���3��(�i�T��� x���ï���ү��  �A�,�e�P�����~� �����ƿؿ��=� (�a�s�VϗςϻϞ� ������� �9�K�.� o�Zߓ�v߈��ߴ��� ���#��G�2�k�N� `������������ �
�C�&�8�y�d��� ������������ć�DBGDEF �|$�:!"�$6 _L?DXDISAQ�#���#MEMO_AP�K�E ?$�
 H�������"ˀISCW 1}$�%�� oy�M�����QE_MSTR �~�m%SCD 1���T/�x/ c/�/�/�/�/�/�/�/ ??>?)?b?M?r?�? �?�?�?�?�?O�?(O O%O^OIO�OmO�O�O �O�O�O _�O$__H_ 3_l_W_�_{_�_�_�_ �_�_o�_2ooBoho So�owo�o�o�o�o�o �o�o.R=va ����������<�'�`��MJPTCFG 1�+�]�%�����MI/R 1�%Ԁp�@T�q���T��< G ?� �%��t�7�q�� i������������� 1�C�֟��j�L�V�x� ��P�����ί��0� T�E �q����8��� ������򿐿����  �B�p�R��ϵ���Z� |���п����6���>� l�R�d߆߈ߖ����� �ߞ���2���@�z� `����������� +�=��������X�b� t�������������* ��o�6��� ������
 @nP���Xz ����4/�,/j/@P/b/�/�/���K��;���  �/���LTARM_�"�̅� �"����6?�>4��METPU ; T����%���NDSP_ADC�OLX5� c>CMN�Ty? l5MST ��-�?���!�?|�4l5POSCF�7=�>PRPM�?�9[STw01���4܁<#�
gA[�gEwO �GcO�O�O�O�O�O�O _�O_G_)_;_}___�q_�_�_�_�_�Ql1S�ING_CHK � |?$MODA�Q3����#5v�eE{�&bDEV �	��	MC:>WlHSIZEX0�-��#eTASK �%��%$1234?56789 �o�e�!gTRI����� l̅%&�0O2}���cYP�a���9d"cEM_IN�F 1�7;a�`)AT&FVg0E0X�})�q�E0V1&A3&�B1&D2&S0�&C1S0=�})�ATZ�#�
�H@'�O��qCw��A�@��b�ˏ���� � &�������3��� ۏȟڟ������"�4� �X�����A�S�e� ֯៛��C�0���� f�!���q�����s�� ������ͯ>��bϙ� sϘ�K���w������� �ɿۿL����#ϔ� ��Y�����ߩ߳�$� ��H�/�l�~�1ߢ�U� g�yߋ���� �2�i� V�	�z�5���������~�.ONITOR�0�G ?kk   	EXEC1�2�2345��`789���( �4�@�L�X��d�p�|�2��2�2�2�2��2�2�2�2��2�3�3�3�(#aR_GRP_�SV 1��{ �(�Q�4����Ҿ�~?���E?��\��3�+���a_Ds�n~�ION_DB-`��1m�1  �� �Fh"$ �++e��0Fh��N �8�2)Fi-ud1�}e�/�/�/1PL_NAME !�e�� �!Def�ault Per�sonality� (from FsD)b"P0RR2�� 1�L68L�@P�!?`
 d�2-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�Of#2)?�O�O�O__@,_>_P_b_t_f"<�O �_�_�_�_�_�_
oo�.o@oRodotl�" D�_�n
�o�of$P�o �o $6HZl ~������� �o�o2�D�V�h�z��� ����ԏ���
�� .�@��!�v������� ��П�����*�<� N�`�r�����e�F���ïխf"d�� ������(�6������ �m���j���V� ������Ŀֿ������:Ϸ�]�m�f"��	`���ϲ��σ�:�oAb)������c' A� � /�	23��)X ����E ���X, �@D�  t�?��z�n�?f |�f!AI��t�j��;�	�l��	 �� � �h�Y !0����� � x � �� ��ҷK_�K }K7X��K��J��?J�+Ƀ�%���ԯC�@�6@��
�\��(E@��Sє��.��=�N��������T;f�a������$��* � ´  �1�>�����z�w����<�
��� ��!�/���1�yD� � �  � W �`�#H �l�����-�	'� �� ��I� ��  �0�&�:��È��È=�s����0�@��@��%�f���f�(��2�+�a!v  '��Y��@!�p@����@��@��@���C��C� �W� C��C��C��=f �A�����'��9"T�Bb $`/��Lf!Dz�� o��~������h���A �кD��  X ,f �?��ffG�*/</� !}�q/�+1�8~`�/�*>��$��(�	(~`�%P�(�������>�$���W�<��	<S�;���9<��<#*o<��M,3@�K;|��f��"�,�?fff? ?y&�0T�@�.�2�J<?N\��5 5	��1��(�|��?z� �?j7��[/0OOTO?O xOcO�O�O�O�O�O�O{h�5F���O2_�O V_�?w_�9I_�_E_�_ �_�_�_oooLo7o po[o�oo�o�oU�o �o��m_3�_Z�o~0���O*��& Q/�wl��q
�m.��+�d�V���Aa0��5�uCP���L�č?����#��Y[�/Ӄ6�B]�D��CC3� z����y�����@I�l�����A��A���PA �R?�1>�-8������ÍO\����Q�����#�
�؞���AиR�A���C;����Q섟"\�)C0����qBo
=��Q�����8�Hp���G� H��0�H��E1� C�&�Hy���I��H���%F�� E,��s�]�i�EI���@H���H���E# D� 7�د�կ���2�� V�A�z�e�w�����Կ �������@�R�=� v�aϚυϾϩ����� ����<�'�`�K߄� oߨߺߥ�������� &��J�5�G��k�� ����������"�� F�1�j�U���y����� ��������0T ?x�u�������P�(��3�(��	4��<�<�̷�t�Ӂ3�� ����ʭ��Ӂ� �&n�
/4�f4yϱ$-$)d/R/��/v/�/�,ՅPD2P�.�a�o?Z?=?(?a?L<?g?n?�?�?��?�?�?  �����?�?+OOOO:OsO@?�o�O�O�O�L7�O��O_�O _F_4_JQ�L_^_�_�_�_�_�_��Z  2jOo  QB��}���Cq���Ӏ@��RoӀMqko}o�o^o�oҌo�o�o�/Aӄ�TRӀӀ�aӀ؎
 I���� ����)�;�M�_�pq����sq ����1��"�$MS�KCFMAP  �$%� ��Vsqoq莼�ON�REL  �%�Ӂ�P��EXCFENB�
у����FNy�'��JOG_OVLIM�d���d��KEY�zq�z�_PAN��������RUNa����SFSPDTY�� '����SIGN|��T1MOTc�����_CE_G�RP 1�$%Ӄ\dOh�\O�����T ��ɯ�����#�گ G���<�}�4�����j� ׿�����Ŀ1��*� g�ϋϝτ���x����������f��QZ_�EDIT�͇��T�COM_CFG 1�ɍ~vv߈ߚ�}
V�_ARC_"���%P�T_MN_oMODE��0�UAP_CPL���4�NOCHECK� ?ɋ  �%�3�E�W�i�{�� ��������������/�A��NO_WA�IT_L�K�6�N�T^��ɋu|��_7ERR@�2�ɉ�Q� ������a��4F��MO������|t5�!�������"��B�o-B�^�/����<���?�l�Knp����_PARAM��ɋ�/�2t8��_^ =�P345?678901x� �s����//`�9/K/'+t7�}/��,"�/��ODRD�SP���0�OFFSET_CARAМ��&DIS�/�#S;_A��ARK�L��OPEN_FIL�E0h���Lִ�OPTION_IO�����m0M_PRG ;%Ɋ%$*�?�>�I3WO50�F��0� �5���2���0@�'A	 a���C���#�� �RG_DSBL  Ʌ�v|rO�!RIENTTO��!C�mpҁ,a� �UT_SIM_D�u7Ђ��� V� LCT ���H��4����I�%y��A_PEqX��?TRAT��� d0�T� UP� ��N�pK���i_{_XrfS`�gq�2�m�}]�$�2?���L68L@P>�C
 d�/�_ oo*o<oNo`oro�o �o�o�o�o�o�o &8J\��2�_� ������
�� .��{X�j�|����� ��ď֏������πH�X��PX�~��"P k�����̟ޟ��� &�8�J�\�n������� ����������"�4� F�X�j�|�������Ŀ ֿ���ɯۯ0�B�T� f�xϊϜϮ������� ����,�>���EC�}ߏ�SI�� �ޤ�����b�bݢ/3��W�
�@L�v�l� ~��������J�Q0�'�)L�	``�Z�xl�~���:�o�A���������KA��  ���T�POOP1��[�v���TH��E�=DX,? @D�  2�4�,?�D442�9�h;�	l�	�@� � �h�_`� ��� � x? � � ��J�H�H2�-�HL��H�l�H�WG����=�3Ho��JC�R�@p�@ז@�PT1���0@�S �>PP%ICUB��<��K�`�@��a�y��  �  _�  � #�0��*&�H/�	'�� � f"I� �  ����=��͊/�+�@�/� �>A�/DM+>B���N�@4?  'x0L4�0}C�@C�� C�C�C�Y?k?D� � �A�!�������/��B�@�1 �����!
ENz�-O �QO<OaO�O^/p(�1<�E�S� �<��1��P.   �?�faf��O�O�O 7��/_A[sA8�W_eZ>��' �FjJ(��UP�X�I�����#�T[��<��	<S�;��9<��<#*�o<��5�\@�	k:��#�R���?fff?� ?&�D`�@�.Vb�?J<?N\�be:� �2?aKjI:�o8�o (g~_�o�o�o6 !ZE~�{�� �����o�o�o� h����w�����ԏ�� я
���.��R�=�v� a�?��o�e+��O�����<�N�`�r�Z���@_��l� /�ȯ�+��ׯ�"����A`>��?�C�s�
�<П��?�ء�����̿n	�/X�j��B�D90CC��ޚ�������^�@I��*����A���A��PA ��R?�1>��-���������O\����Q����#�
�����A�иRA���C;���Q�B���0\)C0����qBo
=���Q�������Hp��G�� H�0�H��E1� C����Hy��I���H��%F�� �E,�1߯i�E�I��@H����H��E# D����ߨߓ��� ���������8�#�5� n�Y��}������� �����4��X�C�|� g��������������� 	B-fxc� ������ >)bM�q�� ���/�(//L/ 7/p/[/m/�/�/�/�/ �/�/?�/6?H?3?l? W?�?{?�?�?�?�?�?tO��(��3�([���T��BE�5�̷�2ODOX�3���8^OpO~B�ʭ�O�O�X�� &n�O�O4�f4yϱ�M �I"__F_4_j_X\��%PbP�^�����_@O�_�_�_o
l?%o�,oeoPouo�o�o  ���ʞo�o�o�o �o1�_��dR�v|7����������
��R�@�pv�d�����  2(�я  BG�;�G�C/�D�X�@K��"�@4�F�X�j�{����������ɟ۟���X�J��X�X���X���
 �W�i� {�������ïկ������/�A���1� ����K1��"�$�PARAM_ME�NU ?�E��  �MNUTOOL�NUM[1]݆���F~������AWEPCR��.�$INCH_RA�TE��SHEL�L_CFG.$J�OB_BAS߰ �WVWPR.�$CENTER_�RI������AZI�MUTH OPT�B����ELEV�ATION TCگ���DW�TY�PE SN�AR�CLINK_AT~ �STATUSǳ~]�__VALU߱�̰LEP��.$WP_�����U�̢� �����������7�2��D�V��z�SSREL_ID  �E��Q���USE_P�ROG %��%x{��ߏ�CCRT����Q����_HOST7 !��!��5���T�P��Q��*��S����_TIMEsOU�Ս�  z�?GDEBUG�Љ����GINP_FLgMSK����TR����PGd�  ����$�CH����Q���z�tߪ����� ����(:c^ p�������  ;6HZ�~ ������//� /2/[/��WORD� ?	��
 	�RS�CPN<n�BMAIW��#3SU&��#TEt�C�STYL C�OL0eW(�/W�TR�ACECTL 1��E�� �P ��6DT �Q��ED0!0D� � �S���QQ6�[<�f�Qy01�q? �?�?�?Q5�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c�u��� ������Ϗ�����)�;�M�_�q�S36L�EW���5��3 � �6_UP ��<;b������ #���&�0�M$a���R�\0R�  ���)_DEFSPoD ���2��o  �z�INؐ?TRL ���a��8!�h�PE_CO�NFIܐ�7����M!b,LID�ٓ���	ĨGRP� 1�9 �lM!A>ff���\�
=D��  DZ� DZ
�@�
�M d!�0?�O�������H�8"�$�i� ´����m�B��̱��������̿��&�B3�4�$�]�o�Y� <<j��tϭ�pϪ� ������ό��O��_߅�p��z�ӳ�M 
���ߊ������5�  �Y�D�}�h����@���������*�)<��
V7.10b�eta1�� �A�k�\�B
�y�(�Y�?&ffp�/>.{X�
������X�B!�~��A{33A�&�(�h� -���������*��pM"��3�EWM$ғ�KNO?W_M  0�薾ȤSV �:�%����� ��IM"G��UM�=�(�	��?���.��* ����&M#�)�Y�@)����M % .ѐȡMR�=�$����f/�x+��ST�1 15�<9^ 4�( )�o��/�/�/
?�/? !?S?E?W?�?{?�?�? �?�?O�?�?>OO/O tOSOeOwO�'2�,��/���<�O�O� A3�O�O�O�O�'4_-_?_Q_�'5n_�_�_�_�'6�_�_�_�_�'A7o&o8oJo�'8gopyo�o�o�'MAD��� ȕ�EOVLD  ���P}�$�PARNUM  ��+?Q�#SCHy ȕ
�wlq�y��uUPDl=u�|��E_CMP_u�����_�'ݥ%�E_R_CHK3�ۣ0 �G�0�B�RSA ��ȡ_MOp����_����E_RES_G
� ���
��p�"�� F�9�j�]�o�����ğ ���۟����o��@���1��PN�m� r��mP��������P ̯���`�*�/� �f`J�i�n�惹`��x�����V 1���|ށ�@]s8��THR_INRA ��q]مd�MASmS)� Z=�MN(��[�MON_QUEUE �����Ъ!ބN*�Un�N8kƔȫ�END��Ώ���EXE�����pB�E���ϫ�OPTI�O��׋��PROG�RAM %��%���習��TAS�K_It �OCFG ��π�ߵЯDATAx����G2�$�6�H�Z� l�������������� �2���INFOx�혝���� ������������	 -?Qcu���@����N�Z���c ����pK_�ѣ���z�5G��2��D X,	}	x�=��O��@���$� �����0_EDIT �����>��WERFL�����#RGADJ M��AЛ@R$?�]%0�5&��?���?�?���A<��z�%�o�/)(�/s#2�'"	�H��l�!?�8�Aٴ�t$�26*A0/C2 **:L2�??Q3m=2���2�5��+1�9��/�?y=�=�? �?�?�?�?KO�?O5O +O=O�OaOsO�O�O�O #_�O�O___�_9_ K_y_o_�_�_�_�_�_ �_�_goo#oQoGoYo �o}o�o�o�o�o?�o �o)1�Ug� �������	� ��-�?�m�c�u�� ��ُϏ�[���E� ;�M�ǟq��������� 3�ݟ���%���I� [���������ǯ������	�ߖ�𰄿 ����39߿53��ϧ��0�B�o'PREF S�*00
5%?IORITY:��}�9!MPDSP8�'*z��UT��34&�ODUCT����E��&OG_�TG$ �����TO�ENT 1��� (!AF_I�NE��Y�J�!�tcpdߌ�!�ud{ߴ�!iccm���.��XYx#���1)� 0Y1�*�0��S� 6�B��f������ ������!�3��W�>�${���*��x#�)P��/������Y7/�c<��44��(�.A~�",  �u� (}���+%�^��f�x�,9!POR_T_NUM��0��9!_CAR�TREP% �aSoKSTA�� 4�LGSV������#0Unothing�����L�]TEMP �����T��_a_seiban� ,/�</b/M/�/q/�/ �/�/�/�/�/�/(?? L?7?p?[?�??�?�? �?�?�?O�?6O!OZO EOWO�O{O�O�O�O�O �O�O_2__V_A_z_ e_�_�_�_�_�_�_�_|o�VERSI�����M` di�sabled'oS�AVE ���	�2670H78%2J�o�o!$�o�o���o 	x��V��.�eKt���J�c|�o��ܺmb_� 1����`*�p�!�4�F���W�URGE_ENaBЪ�(���WFr�#DO���+�WRГ����WRUP_DELAY �,���R_HOT �%{���#���R_?NORMAL���x�W�&�SEMI6��\���U�QSKIP���#�xo��	o ��(���Y�G�}� ����g�ů��կ��� ��C�1�g�y���Q� ���������	�Ͽ-� �=�c�uχ�Mϫϙ� �����Ϲ��)��M��_�q����$RBT�IF��0RCVT�MOUE�����DCR�Ǿ�� ���6u�C^)C7���@���@�nߒ6悔띶���^��R������-��ÿj���H�3�<��	<S�;���9<��<#?*o<��M�Q 7���y������ ��/�A�S�e�w�������RDIO_T?YPE  ������EFPOS1 +1�ui� xA
 -���G2k�o�* �N����1 �UgN�� �n��/�/Q/ �u//�/4/�/�/j/ |/�/??;?�/_?�/ �??�?�?T?�?x?O �?%O7O�?�?OOjO��O��OS2 1�ԋZO�O_�O6_<�O��3 1��O�O��O,_�_�_�_L_S4 1�c_u_�_�_?o�*oco�_S5 1� �_
ooVo�o�o�ovoS6 1͍o�o�o��oiT�S7 1�"4F���|"��S8 1Ϸ������~���5�SMASK 1����  �� �ՇXNO����)�=�����MO�TE��=�Z�_CFG �a���)����PL_RANG�]��ߛ�OWER ��%�ΐ��SM�_DRYPRG �%%�%^��ԕT?ART �ƞ�UME_PRO����p�=�_EXEC_ENB  ����GSPDI�������Ѣ�TDB����R�Mϯ��IA_OPOTION������.U�MT_݀T��_�2��*�z��9���C�ˀ�����������OBOT__ISOLC"������ֵNAME �%�_���OB�_ORD_NUM� ?Ƙ���H782  ˄h�@h�$�hʬ��h�>�PC_TIM�E�ם�x��S23�2z�1����L�TEACH PENDAN��v�A��~�]�H@Ma�intenanc�e Cons˂���ˆ"�DDNo Use~�E��i��{ߍߟ߱ߵ���NPQO#���A�!���oCH_LL��U�樀	3���!U�D1:Y� �R܀VgAILI���žU�SR  %������R_INoTVAL����������V_DAT�A_GRP 2�X%���X�D��P�� W���{�f�%������� ��������$& 8n\����� ���4"XF |j������ �//B/0/R/x/f/ �/�/�/�/�/�/�/�/ ?>?,?b?P?�?t?�? �?�?�?�?O�?(OO LO:O\O^OpO�O�O�O �O�O�O_ _"_H_6_�l_U��$SAF_DO_PULS���V���X��Q�PCANd������SC���(�}���ˀq����x�C�C��˂ p�o0oBoTo foxoo�o�o�o�o�o,�o�����be�$!r �dt:ql�(s�� @��fx�Ȝ~Ny� D�t_�_ @�T������T D��*�S�e�w��� ������я����� +�=�O�a�s�����`u/2���ǟ�і��C���;�o�2���p����
�?t��Di���a�C��  � � ��Cђax��Qa�s��� ������ͯ߯��� '�9�K�]�o������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��π��������1�2�� aZ�l�~ߐߢߴ��� ����9�u�(�:�L� ^�p��������2�0�D��N�	�� -�?�Q�c�u������� ��������); M_q����� ��%7I[ m�����D� �/!/3/E/W/i/{/ �/�/
��/�/�/�/? ?/?A?S?������r �?�?�?�?�?�?�?O #O5OGOYOgIzO�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo`o5�艟9�ko�o�o �o�o�o&8J \n�����pj��o��2����S����	12�345678+��h!B!ܺ�4���`��|��� ����ď֏����� �o5�G�Y�k�}����� ��şן�����1� C�U�f�$��������� ѯ�����+�=�O� a�s�������h�z�߿ ���'�9�K�]�o� �ϓϥϷ��������� ��#�5�G�Y�k�}ߏ� �߳����������� 1�C�U��y���� ��������	��-�?� Q�c�u�������j��� ����);M_ q������� ��%7I[m �������/ !/3/E/W/{/�/�/ �/�/�/�/�/??/? A?S?e?w?�?�?�?�sm��?�?q/OO�*OF�Cz  B}pqj   ��hu2�bm�} ph�
�G�  	��r2�?�O�O�O�OokK>�_Dlo�<��O B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o'_�o�o�o �o(:L^p ������� ��$�>ISB�1�AiB�<S��$SCR�_GRP 1���8� � �� �SA �dE	 ��������� �1B���SG��ۏɏ�N:M�s@��D^@�D/^��E��� \�ARC Mat�e 100iD/�1450ҁAM��ҁMD45 �678SC
12�345��9��Ӆ E����KyBד_��SF �߃� S��Ó��Ӂ�	yJ6�H�Z�l�~�~SD��H���������Əǯ���Ά�oSAگC�֯�g�N���v�B�M@Ɛ����ɴ��A^@ؿ c @S@𵬁@��F� ?PŬ�HM@�)�ۺ��F@ F�`S�[�~��jϣ� �ϳ���������!ߤ��� �L�7�I�[�m�B�{���߬�����	� ���?�*�c�N��r� ��_��)������dGA�@��0�SB�@PG7H�_�!�@�4p�M@Ȇ�����߃�?��SDA�����$���� QƒSAA 3E��!h�t�U (�  ������ �$�SF_�EL_DEFAULT  锿��S@~@HOTSTRL�#^�EMIPOWERFL  BExX?�WFDOM� �RVENT? 1�����w� L!DUM�_EIP.���j�!AF_INExL/SD!FT��@./d/!���/ ��S/�/!RP?C_MAIN�/�(q��/�/�#VIS�/�)��/H?!TP&;0PU??�d7?�?�!
PMON_POROXY�?�e�?��?[2�?�f�?,O!�RDM_SRV�-O�gOxO!RȲ��O�hgO�O!
�� M�?�i�O_!RLSYNC_���8�O\_!R3OS��\�4K_�_�!
CE]0MTC�OM�_�k�_�_!=	�RCONS�_��l�_@o!�RWA'SRCGO�m/o�o;!�RUSB�o�n{o�ow/�o;C�o�o %Jn5�Y��:RVICE_K�L ?%� (�%SVCPRG1����u2�
��p3-�2��p4U�Z��p5}����p6�����p�7͏ҏ�p����9�"��t�OJ��q� r��q����qG��q o���q����q��:� �q�b��q����q7� ���`�گ����� ��*��؟R�� �z� �(����P�ʿ�x� ������ȯB�D� ���r�p��p���� <��������	�B�-� f�Qߊߜ߇��߫��� �����,��>�b�M� ��q��������� ��(��L�7�p�[��� ������������� 6!ZlW�{� �����2�V�z_DEV ���MC:���T4��pGRP 2�����p�bx 	� 
 ,�^��� �/�&///\/C/ �/g/�/�/�/�/�/�/ ?�/4??X?j?��? E?�?�?�?�?�?OO OBO)OfOMO_O�O�O �O�O�O�O�O_q?_ P__t_[_�_�_�_�_ �_�_o�_(ooLo^o Eo�oio�o�o�o�o3_  �o6ZAS �w������ �2�D�+�h�O����� �oy����ߏ�� @�R�9�v�]������� П����۟�*��N� ��C���;�����̯ޯ ů��&�8��\�C� ����y�����ڿ��ӿ �g�4�F�-�j�Qώ� uχ��ϫ������� �B�)�f�x�_ߜ߃� ����)��߭��,�� P�7�t��m����� �������(��L�^� E�����w���o�����  ��6ZlS �w�����p�D��d Ԗ�	2{f������O%��/�����4!�4%D/R' </r/`/�/�/�/�)/ �/0)�/??>?,?N? P?b?�?�/�?�/�?�? �?OO:O(OJO�?�? �O�?pO�O�O�O�O_  _6_xO]_�O&_�_"_ �_�_�_�_�_oP_5o t_�_hoVo�ozo�o�o �o�o(oLo�o@. dR�v�� � $���<�*�`�N� �������t���p�ޏ ��8�&�\����� L�����Ɵȟڟ��� 4�v�[���$���|��� ��¯į֯�N�3�r� ��f�T���x������� �:��J��>�,�b� Pφ�tϪ����Ϛ� ߖ��:�(�^�L߂� �ϩ���r����� ��� �6�$�Z�߁���J� ������������2� t�Y���"���z����� ������:�1��
 ��R�v��� �6�*:<N �r����/ �&//6/8/J/�/� �/�p/�/�/�/�/"? ?2?�/�/?�/X?�? �?�?�?�?�?O`?EO �?OxO
O�O�O�O�O �O�O8O_\O�OP_>_ t_b_�_�_�_�__�_ 4_�_(ooLo:opo^o �o�o�_�oo�o �o $H6l�o�� \~X��� �� D��k��4������� ������^�C��� �v�d����������� ��6��Z��N�<�r� `���������"��2� ̯&��J�8�n�\��� ԯ�������~���"� �F�4�jϬ���пZ� �ϲ���������B� ��iߨ�2ߜߊ��߮� �������\�A��
� t�b�������"� ��������:�p�^� �������������  "$6lZ��� �������  2h���X� ���
/�/p� g/�@/�/�/�/�/�/ �/?H/-?l/�/`?�/ p?�?�?�?�?�? ?O D?�?8O&O\OJOlO�O �O�O�?�OO�O_�O 4_"_X_F_h_�_�O�_ �O~_�_�_o�_0oo To�_{o�oDofo@o�o �o�o�o,noS�o �t����� �F+�j�^�L��� p�������܏��B� ̏6�$�Z�H�~�l��� �
�۟������2�  �V�D�z�������j� ԯf��
���.��R� ��y���B�����п�� ����*�l�Qϐ�� ��rϨϖ��Ϻ���� D�)�h���\�J߀�n� �ߒ���
������� ��"�X�F�|�j���� ��������
��� T�B�x������h��� ������P�� w��@����� �X~O�(� p�����0/ T�H/�X/~/l/�/ �/�//�/,/�/ ?? D?2?T?z?h?�?�/�? ?�?�?�?O
O@O.O POvO�?�O�?fO�O�O �O�O__<_~Oc_u_ ,_N_(_�_�_�_�_�_ oV_;oz_ono\o~o �o�o�o�o�o.oRo �oF4jXz|� ��*���B� 0�f�T�v���Ï� �������>�,�b� ����ȏR���N�̟� ����:�|�a���*� ��������ȯ�ܯ� T�9�x��l�Z���~� ����Ŀ�,��P�ڿ D�2�h�Vό�zϰ�� ���Ϡ��Ϝ�
�@�.� d�R߈��ϯ���x��� �������<�*�`�� ����P��������� ���8�z�_���(��� ������������@�f� 7v�jX�|� ���<�0� @fT�x��� �/�,//</b/ P/�/��/�v/�/�/ ?�/(??8?^?�/�? �/N?�?�?�?�? O�? $Of?KO]OO6OO~O �O�O�O�O�O>O#_bO �OV_D_f_h_z_�_�_ �__�_:_�_.ooRo @obodovo�o�_�oo �o�o*N<^ �o�o��o���� �&��J��q��:� ��6���ڏȏ���"� d�I����|�j����� ��֟ğ��<�!�`�� T�B�x�f�������ү ���8�¯,��P�>� t�b���گ��ѿ���� ���(��L�:�pϲ� ��ֿ`��ϸ������� $��Hߊ�o߮�8ߢ� ���ߴ������� �b� G���z�h����� ����(�N��^���R� @�v�d������� ��� $�����(N<r `��������� $J8n�� �^����/�  /F/�m/�6/�/�/ �/�/�/�/?N/3?E? �/?�/f?�?�?�?�?��?&?OJ?L1�$S�ERV_MAILW  T5J@�0H�OUTPUT?H�0HRV �2��6  M@ �(�1O�O4DTOP�10 2�I d P?�O�O__ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9K] o�������5ιEYPE`LNEFZ�N_CFG ��5MCL4oB�?GRP 2�%��� ,B   A�e�L1D;� B�f��  B4L3�RB21�FHELL���5��@�O<�ΏK%RSRݏޏ��)��M� 8�q�\�������˟����ڟ���7�I�[��  �+�[���X��i��� L0��PŢơL8q�2L0d��������HK 1��� ˯@�J�D� n���������߿ڿ� ��'�"�4�F�o�j�|���ϊ�OMM �����Ϗ�FTOV_�ENB?D�A��O�W_REG_UI���2BIMIOFW�DL�����h�3�WAIT����oE^��Z@��DX�TIMn�����VA>@|i�3�_UNIT������LC�TRY���4@MON�_ALIAS ?5e���@heOM� _�q��J;������ ���� �2�D�V�� z���������m����� 
.��Rdv� 3������ *<N`��� ��w�//&/8/ �\/n/�/�/=/�/�/ �/�/�/�/"?4?F?X? j??�?�?�?�?�?�? �?OO0O�?AOfOxO �O�OGO�O�O�O�O_ �O,_>_P_b_t__�_ �_�_�_�_�_oo(o :o�_^opo�o�o�oQo �o�o�o �o6H Zl~)���� ��� �2�D��h� z�������[�ԏ��� 
��Ǐ@�R�d�v��� 3�����П⟍��� *�<�N���r������� ��e�ޯ���&�ѯ J�\�n���+�����ȿ ڿ쿗��"�4�F�X� �|ώϠϲ���o��� ����0���T�f�x� ��5߮��������ߡ���,�>�P�b���$�SMON_DEF�PROG &������� &*SYST�EM*i�����<{�RECA�LL ?}�� �( �}3xco�py fr:\*�.* virt:�\tmpback���=>192.1�68.56.1:?13648 � �X2�D��}4��a������������ }�8��s:orde�rfil.dat�v�����/AS}/��mdb:s�� ���`���z�� �.@Re���� �������~�*/ </N/as/��/�/ �/�r�&?8?J? ]o ?��?�?�?� �v//"O4OFOY/k/ O�/�O�O�O�/�/|? ?�O0_B_�Og?�O
_ _�_�_�_�?�?�O�O ,o>oPocO�_�Oo�o �o�o�Ot_�__(: L__�o�_��� �_�_xoo$�6�H�[o mo��o����Ə�o�o ~ �2�D�Wi�� ����U����� ��.�@�R�e� ���� ����Я�v����*� <�N�a��������� ̿ߟ�z��&�8�J� ]�o�
ϓ��϶���ۯ ���"�4�F�Y�k� �Ϗ��߲���׿��� �ߟ�0�B���g��� ��������x߅�� ,�>�P�c�����ߪ� ��������|��(: L_�s����� ������$6H[� m����������� t� /2/D/Wi/��/�/�/U.�$S�NPX_ASG �2�����!��  0��%��/?  ?���&PARAM ���%�! ��		;P����o4�� OFT�_KB_CFG � ��%�#OPI�N_SIM  
�+j2�?�?�?�3�� RVNORDY?_DO  t5�5�BQSTP_D�SB�>j2HO�+S�R ��) �� &n:�O��&T�OP_ON_ER�RO�FPTN ��%�@�C��BRING_PR�M�O#BVCNT_�GP 2��%l1 0x 	DO?_�-_�f_Q_�_�'VDPROP 1�C9m0{Q �1m_�_�_�_�_o4o 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu����� ����)�;�M�_� ����������ˏݏ� ��%�L�I�[�m�� ������ǟٟ��� !�3�E�W�i�{����� ��دկ�����/� A�S�e�w��������� ѿ�����+�=�d� a�sυϗϩϻ����� ���*�'�9�K�]�o� �ߓߥ߷��������� �#�5�G�Y�k�}�� ������������� 1�C�U�|�y������� ��������	B?�Qcu���RPRG_COUNT�6s��B�	ENB�O��M��4�_UP�D 1�nKT  
��ASe� �������/ /+/=/f/a/s/�/�/ �/�/�/�/�/??>? 9?K?]?�?�?�?�?�? �?�?�?OO#O5O^O YOkO}O�O�O�O�O�O �O�O_6_1_C_U_~_ y_�_�_�_�_�_�_o 	oo-oVoQocouo�o �o�o�o�o�o�o. );Mvq��� ������%�N� I�[�m���������ޏ�ُ돷_INFOg 1�/ �� �R�=�v�a�������!�������"�B�o-�B�^������YSDEBUG�� 0���d��S�P_PASS��B?�LOG ��/9  r�����  ����UD1:\x���_MPC$��/����/[�Я �/��SAV ��'����G�_����f�SVԛTEM_TIME 1�'�]: 0� �����үr�4�SKM�EM  /�.G�  ��%s���\Ͽ��� @����h������"��P׿
A���;��D�V�*��nʟ�����ϐ�ϸ���^��E�� W�������+�=� O�a�s߅ߗߩ߻����������{�9�K� ]�o��������� �����#�5�G�Y�k��}���T1SVGgUNS*�'����ASK_OPTION� /���_DI�����BC2_GRP �2�/�Q�%��@�`�C�:��BCC�FG �� 9����`��� �����!E 0iT�x��� ��/�///?/e/ P/�/t/�/�/�/�/�/ ?��,!?�/T?f?�/ C?�?�?�?�?�?׮O ���0O2O OVODOzO hO�O�O�O�O�O�O�O _
_@_._d_R_t_�_ �_�_�_�_�_o�_o o*o`oFh10to�o�o �o�oFo�o�o�o" FXj8�|�� �����0��T� B�x�f�������ҏ�� �����>�,�N�P� b�������roԟ�� �(���L�:�\���p� ����ʯ���ܯ� � 6�$�F�H�Z���~��� ��ؿƿ����2� � V�D�z�hϞόϮϰ� �������ҟ4�F�d� v߈�߬ߚ߼����� ��*���N�<�r�`� ����������� �8�&�\�J�l����� ������������ "XF|2ߔ�� ��f�B0 fx�X���� ��///P/>/t/ b/�/�/�/�/�/�/�/ ??:?(?^?L?n?p? �?�?�?�?��?O$O 6OHO�?lOZO|O�O�O �O�O�O�O_�O2_ _ V_D_f_h_z_�_�_�_ �_�_�_o
o,oRo@o vodo�o�o�o�o�o�o �o<�?Tf� ��&����� &�8�J��n�\����� ����Əȏڏ���4� "�X�F�|�j������� ֟ğ�����.�0� B�x�f���R��Ư� �����,��<�b�P����p���A��*S�YSTEM*��V9.0055 ���1/31/201�7 A v  ���K�TBCS�G_GRP_T �  \ $E�NABLE�$�APPRC_SC�L   
$�OPEN�CLO�SE�S_MIN;F2'�ACC���PARAM� ����MC_MAXo_TRQ�$dį_MGNk�C�A�Vw�STALw�B{RKw�NOLDw��SHORTMO_GLIM�ʧ�h�J�����PL1��6���3���4��5��6��7���8k�����O� $D�E�E���T��b�PATH�^�w�m�w�_RAT�IOk�s�T� 2 	$CNT�aA�����m�INXѯ_UCA���C�AT_UM��YC_ID 	����_E����6����~��PAYLOA���J2L_UPR_7ANG6�LWA�?��3�O�x�R_F2LoSHRTv�LOD����}��Ӌ���ACRL_S�ؽ���+�k�wHVA�$Hx�^��FLEX�BѻJ2� P�B�_F��$��_F�TM��&��$?RESERV�>��;������� :$��LE1N.�z�;�DE|����;�Yғؔ��SLO�W_AXI��$�F1��I��2��1�������MOVE_�TIM��_INE�RTI��
�	$D~TORQUEX��3��#I��ACE�MN��%E�%Ep	V��d�A�R�TCV��Rt��(��
��T@�RBJ���	M���,��J_MOD8����� dR�y�2��PpE����\�X��AW�gQJK@��mK��VK�VK�gJJ0���JJ��JJ�AA��AAf�AA%�AA �t�N1�N �d�#���E_NU�����CFG� �� $GROU�Pc�SK��B_C�ON�C��B_R?EQUIRE����BU��UPDAT�T�EL}  ��%� $TJڧ�� JE��CTYR��
TN F�&��'HAND_VB���OP� �$oF2x�3�m�C?OMP_SW��@��R�� $$Ma�e�R�Î8���<� ��5�¼6A_.�h�DT�<q�A��A��A��QA���0��D��D��5D��P��GR�ǂACST�ǂA�ɂAN��DY���x��4�5A� ��s��s��2�B��R����P���Հ� �)�2�;�h��c �0i�\� 7x�U6��QASYM��
�TС��мݎ���_SH�"�����̀�TU8����%�7�J�>���P�pcfio�_�VI83�h6þ`V_UNI���d�{�JU�bU�b���d�� �d v����������su��� �A��H7R_T��	N2�qL���DI����O�t8K¢p�#
  �2I�QAz����q �S��s � B� �p � � f1MEBe���pr�QT�pPT&`r a�>���~$A�5`C�^�R�T4`�! $DUM�MY1�$PS�_ RF��$�����FLA� Y�P_��F�$GLB_T�0�u΅>���pB�; 1�q X��'�STf� S�BRv�M21_V�T$SV_ERba�O(`�,�CL���Ap O�r�pGL��`EW� 4 �$H�$Y�2ZB�2Ww��x�b3A����e�Y�U]� �oN��)`$GI�0}$]� �� Y���� L�h���'b}$F'bE^��NEAR_ N��yF�\ TANC�Ҟr��JOG���� ��� $JOI�NT�&  W�MwSET�  ��E�� S��qϑ|� ��  �Ue?�� LOC�K_FO��m1�pB�GLV3GL��T?EST_XM�j�'EMP=�Ϣ悎��$UC�\���2� ������i0�����CE| Ó�_ $KAR�M�sTPDRA`�3�*��VEC~�D�.�IU����!CHE��TO�OL��i�V��RENK�IS3;���6�N��ACHP���v�1O��F���29����I��  @$R�AIL_BOXEz�� ROBOƤ�?��HOWWA�R��屖���ROLM���q!��¡!Ӱ���J�O_F� !k �rG�CHK�]6� �RN�Oo�!W���?�C��sZ�KOUR�����Q��"�!��$PIPǦN]�Ӳ�� ���V�@�CORDEDH����u�6�p� O�p  D ̀OBA�#�������p̀��'`�!SYS���ADR�!�p>�TC}H�0  ,oSEN�r#�A��_���d�z!�!y�VWV�A� � �9�]��uPREV_�RTA$EDI}T��VSHWR�!��&��]q��`D�(�.Q��6Q$H�EAD8amp��Ha��KEq�|�CPS�PD�JMP�Ld�u�Ra �t��T�\�IРS�"C20�NEr��!�'TIC�K���QM�!%�8�H=N�� @�W�~%�_GP��ʶ$�gSTY^ү�LO��:��� t 5
��Gj�%$�Ѳ�u=��S�!$�a Jp-����p��P�P��SQU-������aTGERCB��1� S�$ ����']�'-`�>pOC�6�bP�IZ��������P�R������S��PU��a��_DO�c�XuSN�K�vAXI��/���UR� p�" 찕�"�]1� _`�4ҋET5P��ЦU���F�W��A�A�Q���ĳ��!&�T{SRE4lu� �9��:��6�	�2� �7��9��9�G� G�'F"TIF �R&��4CE op2oDoVds1SSCЀ�  h� DS���4���SP�p"%A	T@�2���c⅂�ADDRESs�B���SHIF�#�_W2CH� �It!�TU�I�1 �W�CUSTOTVs1V��I�r U���6!��P
Ϫ� �"�����! \����� ���,��!�2CSC���Y�*��2�1�TX_SCREE��"�p=�TINAO����T4��r Fj�Q9_6"vP# TI�/� ��4�.���63��4��RRO�@�3а
��1�h�UE?�$# ��PMѧ�SP�4��RSM����UNEaX_�vA�pS_���+F�SA.IIG�S6Cx��B�4 2#�pUErT%�r?�nF��WGMT3pL�a��O@���BBL_r��Wo���& ���j�BO���BLEf"��C밚"�DRIGH��CBRDA�\!CKsGRo�UTEX$ |UQWIDTH�����Ʊ��Jq���UI>�EY6 ��'� dh��Ѐ���Ӱ��BACK�ᡂ�U�E�!�FO���WL[AB�?(!�I����$UR��P���_P'�H�1 ( 	8wq�_��t"�R(�Rq���������f��Q)Om!��)��L�P�U�@7cR���LUqM7cV ERV���D�_PP�fT*��j GE�R�a `�)&�LP�e_E\���)�g��h!�h���iU5�k6�k7�k8�b�Z�6����4����ڎ�S!�)^QUS=R]�+ <��'�1U���#��FO� ��PRIrm��%q�p�TRIPϱm�SUN�p�t,�����p����/��3 -� �-�RSp��G � �T/��u!�rOSF��vR9 �2�so���.f�x������1�	U�a��/$�6�DC�b����sOFFŠ��0���L�O�� 1�.9�����/9�GU.�P���׃��sQ�SUB��H��@SR	T��1���;���sOR��'�RAU� r(�T=�Z��VC� >Ҕ2� ɲ���$���y�8񹳬`C���{�DRIV���@_V�����Ѐ�D~4tMY_UBY3t �����$��19�l0��q	����P_S������BM�A$nb�DEY_�EX�@��3���_MU.�X�An� @USA8��p�[�k0U�xp� �2V�G>gPACINr�!�RG�𦥽�����A���SCp�RE�Rj!o��`���S�3 ^Y�TARGÐP72H���a�R�S�4nP�0`TQ�	o���RmEz�SW��_A���� o���OIq\!A(n v��E$pU�෱�� \Pa�HK��5����W�s��0��sEA��ɷWOR�Pxv����MRCV�AW6 ��`O��M�P�C83	����REF�G(����e�s` cM�Xp�^��^�-�8��Ƶ�_RCʻ���0S!pf�ϓ��~�8����D7 ���gP�TU0 epԕw�OU�����惓 2��2 $U00��Fr�45#�^�K �SULg 5c`CO�0 `6`�]��� �0���Ѫ�a��@q��i�L���$���a���@q�s�?�8|� +5#k� 5#C7ACH2�LOR�&��<�a�A�KQC ��C_oLIMIg#FRj�qTl���$HO�Pz�*�COMM��BO�@��ب �a�F�VP��<���_�����Z����k���WAv{�MP�FAIk�5G��;�AD?�p��IMRE�_���G�P@V�� k�ASY�NBUFk�VRTaD������&SOLo SD_|���WA�P�'ETUO�X�Q�����ECCU�VEM�٠%�k�VIRC�?����B��_DE�LA����p�p�AuG��Rc�XYZM@�5Cc�W3�qsQ T���P�	 
�D9�"�QLASAP�
�� Gl� :�rX�S�a�7�N�_�LEXEE�;�3W�ka5!���FLPIW���F�I����F���PX�9#�<_p�
���8t@s���@ORDB|qȟ��##�� =_0�Z`T�r�B�O|JP6b�VSFE �3>  a0s���c�sUR��@VSM�u#?�rV�R J� f�3�"�5@�r���qLIN��@�W&N�XS屎 A��2���K&SHd`HOL�k(�XVR�tB|��@T_OVRk� �ZABC�C ��"q-1��Zހ�t}D�rDBGLV���Lϒ�R�ZMP�CF�E�0�tL2ޑLN~ ��
� 9Mc��F Ђ`��ɰ4CMCM��C>��CART_Y1���P_2` $	Jw3q4D��}2�2�70`�5`��UX|5�UXEu��6|�5��4�5�1�1�9�1�7A�C�Z�%G �+�$� BYV D.�p H�RRM�{q���HET����P�U'�Q A�I � ��A� P�EAKf���K_ScHI�B��'RV !F�G½B� C�@r2�g1|�����A20��I� S��DXTRAC�E�PV�� -�PH{ER'aJ ,e��THjO|J�$TBC�SG� 2 �����Q�v��� �Q
 ` �_�_�_�_�_�_�_��_.ooRodkwR~S~�\d ��a}?�Q	 HCBdo~�iC  B �R0�o�h�o�kB��o�p��o�jdf  AXp?�w{qW� {������@�@�P:nT�g�z�E�W� �������
����3�	V3.0�0�R	md45N�	*U�M����1�� ��m����  ��֟�wQJ2{c�]6���� � �U�Q ,����E�şp�G�p�����	_� ȯ���ׯ���4�� D�j�U���y�����ֿ �������0��T�?� x�cϜχϬ��Ͻ���@����>�P�X�7� j�|�&ߜ��߬����� 	���-��Q�c�u�� B���������� �U%�7��Q��=�c�Q� ��u������������� ��)M;q_� ������ 7%GI[�� �������// �M/;/]/�/q/�/�/ �/�/�/??%?�/I? 7?m?[?}?�?�?�?�? �?�?�?!OOEO3OiO WOyO�O�O�O�O�O�O _�O__/_e_S_�_ w_�_�_�_�_�_o�_ +ooOo=oso�o//�o �o5/ko�o�o9 'Io]���u �����5�G�Y� k�%���}�������� ׏���1��U�C�e� ��y�����ӟ����� �	��Q�?�u�c��� ������ͯ����o �oA�S���+�q����� ��ݿ˿��%�7�I� [���mϏϑϣ��� �������3�!�W�E� {�iߋߍߟ������� ����A�/�Q�w�e� ������������� �=�+�a�O���s��� ��e���������' K9[]o��� ����#G5 k}��[��� ��//C/1/g/U/ w/y/�/�/�/�/�/	? �/-??=?c?Q?�?u? �?�?�?�?�?�?�?)O OMO_O��wO�O3OaO �O�O�O�O__7_%_ G_m__�_O_�_�_�_ �_�_o!o3oEo�_io Wo�o{o�o�o�o�o�o �o/SAce w������� �)�O�=�s�a����� ����ˏ�O	��-� ׏]�K���o������� ۟ɟ���#�5��Y� G�}�k�����ůׯ�� ����1��U�C�y� g�������ӿ����� �	�?�-�O�Q�cϙ� �Ͻϫ��������� ;�)�_�M߃ߕ�?��� ��i������%��I� 7�m�[�}������������!��E�/� s e�i� i��}�i��$TBJO�P_GRP 2�1�� / ?�i�	�������9� ?� ����+ ��������i�� @e��	 ��CB  ��C�����5GU	i�C� 2BH  A��/��D�,��bB* q��$�7C��  ���c�d�L�i�A �EG+ ��a	���D/�D<Ky/�//#/�/�/��	??�/�/ T?f?%?o?a	�?�?�? �?�?�?�?O)OO!O OO�O[OO�O�O�O�O(�O_g�i�1Q�E	V3.00���md45��*�[P��d�i_tW �G/� G7� �G?h GG8 �GO Gd� �Gz  G�� �G�| G�: �G�� G�� �G�t G�2 �G�� Gݮ �G�l G�* G�� HS�R�F� F@ �F+� FK  �Fj` F� �F�Q � GX� �R�Q^� Gv� G�ĨS�4� G�� G��� G�\ G�� =L��=#�%
]Ae�Js�Yo�kbi�oo�o��E_STPAR�P]����HR�`ABL�E 1	��C`i��h�g ��di�g��hn i�h�p�g	��h
�h�h�ei���h�h�hDa�cRDI�o���o!3EWu�tO��{� ���+��bS��� �z����"�4�F� X�j�|�������ğ֟ �����0�B���Ā ȏ���g��l�~����� N`r���x�bi��NUM  1�U��	 q� C`�D`�b_CFG �
R���@��IM?EBF_TT�a��8���`��VERBc��z����R 1�kO 8f_i�d�2� P���  �� �%�7�I�[�m�ϑ� �ϵ����������!� 3�|�W�i߲ߍߟߵ�������A�����cMD3�E��� k�}��V_I����GINT�����T1�#�5� B��O�a���G_TC������$�P����9�RQ��Դ�_L���@˵�`M�I_CHAN�� �˵ nDBGLV�L��˵�aq ET�HERAD ?*�e� ��`������hq ROUT6��!P�!#A~SNMASK�|˳�255.�GS}��GS�`OOLOFS_DI�P��%�	ORQCTRL ޻7��o-T/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?s</�?�?��?�cPE_DET�AI��PGL_�CONFIG �R�b���/c�ell/$CID?$/grp1�?4O FOXOjO|O2��
�O �O�O�O�O_�O%_7_ I_[_m___�_�_�_ �_�_�_�_�_3oEoWo io{o�oo�o�o�o�o �o�o/ASew �*��������}�O�a�s���@������?я���� ��*�<�N�`���� ������̟ޟm��� &�8�J�\�n������� ��ȯگ�{��"�4� F�X�j���������Ŀ ֿ������0�B�T� f�x�ϜϮ������� �υ��,�>�P�b�t� ��ߪ߼�������� ��(�:�L�^�p��� ��������� ��@��User �View "I}}�1234567890C�U�g�y��������. C����)�2 6���+=Oa����0�3�����@��	h*��4� cu�������5R/)/;/M/_/q/��/��6/�/�/��/??%?�/F?��7 �/?�?�?�?�?�?8?�?��8n?3OEOWOiO�{O�O�?�O�B �lCamera4�*O�O__)_;_M_+�E�Ow_�_�^A���_�_�_�_�_o)  �F���O_oqo�o�o �o�o`_�o�oLo%@7I[m�O��F �	�����%� �oI�[�m�������� Ǐُ돒�wQ��7� I�[�m����8���ǟ ٟ$����!�3�E�W� ���w+k🥯��ɯۯ �����#�5�G���k� }�������ſl��E�) Z��!�3�E�W�i�� �ϟϱ���������� �/�ֿ�wm9��{ߍ� �߱�����|����� h�A�S�e�w���B� �w!I2�������/� A���e�w��������@����������9�� HZl~��I�� ����� 2DV(hz	J	�E0 � ����/�3/E/ W/�{/�/�/�/�/�/ |��@�Ky/.?@?R? d?v?�?//�?�?�?? �?OO*O<ONO�/�E Bk�?�O�O�O�O�O�O �?_*_<_�O`_r_�_ �_�_�_aO��{Q_o o*o<oNo`o_�o�o �o�_�o�o�o& �_�U��or��� ��so���_8� J�\�n�����9�U�� )�ޏ����&�8�� \�n���ˏ����ȟڟ ������U򻕟J�\� n�������K�ȯگ� 7��"�4�F�X�j��  ������� Ͽ����)�;�M�_�   o�w��� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e��w�����������c� � 
�(  �>��( 	 �� ;)_M�q� �����%��� ̹�j| �������/ �Y6/H/Z/�~/�/ �/�/�/�//�/? ? g/D?V?h?z?�?�?�/ �?�?�?-?
OO.O@O ROdO�?�?�O�O�OO �O�O__*_<_�O`_ r_�_�O�_�_�_�_�_ oI_&o8oJo�_no�o �o�o�o�oo!o�o "ioFXj|�� �o���/��0� B�T�f��������� ҏ�����,�s��� b�t���͏����Ο�� ��K�(�:�L���p� ��������ʯ�� � �Y�6�H�Z�l�~��� ׯ�ƿؿ�1�� � 2�D�V�hϯ��Ϟϰ� ��������
��.�u� R�d�v߽Ϛ߬߾���p����;�@ �#�5�G��� ���0frh:\t�pgl\robo�ts\am100�id\arc_m�ate_��_14?50.xml�� ����������0�B�T�E���Y�~����� ���������� 2 D[�Uz���� ���
.@W Qv������ �//*/</SM/r/ �/�/�/�/�/�/�/? ?&?8?O/I?n?�?�? �?�?�?�?�?�?O"O 4OK?EOjO|O�O�O�O �O�O�O�O__0_GO A_f_x_�_�_�_�_�_��_�_oo,o>n`�Ζ� �k�<<w i�?�>k �o>oyo�o�o�o�o�o �o�o5-O}c ���������1�?��$TPGL�_OUTPUT �I�I� a`i�~������� Ə؏���� �2�D� V�h�z�������ԟ@���
��i�a`�6��2345678901A�S�e�w����� ��?�>�ʯܯ� �� $���(�Z�l�~�����:�}��Կ���
�� ��ƿR�d�vψϚϬ� DϺ�������*��� 8�`�r߄ߖߨ�@�R� ������&�8���F� n�����N����� ���"�4�����j�|� ��������\����� 0B��Px�� ��Xj�, >P�^���� �f�//(/:/L/�A�}\a�/�/�/�/�/�/�-@co?#?ij ( 	 &� X?F?|?j?�?�?�?�? �?�?�?OOBO0OfO TO�OxO�O�O�O�O�O _�O,__<_>_P_�_t_�_4��_`xf�_�_ �]�_o*ooNo`o.� �_�o�o=o�o�o�o�o !o%W�oC� �y��3��� �A�S�-�w����q� ��яk������=� ����s���������� ����a�'�9�ӟ%� o�I�[��������� ��ٯ#�5��Y�k�ɯ S�����M�׿�ÿ� �}��U�g�ϋϝ� wω���1�C�	�ߵ� '�Q�+�=߇ߙ��ϝ� ��i߻�����;�M� ��5���o����� ���_���7�I���m� �Y������%����� ��3i{�� ��K�����/�R�$TPOF?F_LIM �P�>�Q��J�N_SVN  ��$`P_MON7 �Ub���2�%JSTRTCHK �U�`/hVTCO�MPATu�dVWVAR ��"(y � �:/Y�J_D�EFPROG �%�%MAI�nOLDADUR�AQ/�_DISP�LAYU�j"IN�ST_MSK  �, �*INU�SER��$LCK��,�+QUICKM�EN"?�$SCRE�A0�U "tpsc�$�!\0a9`�r0_v9ST�`R�ACE_CFG ��"$Y	�C$
?��8HNL� 2y*�P�1)+  O"O'O9OKO]OoO�O��O�J�5ITEM �2K �%$�12345678�90�O�E  =<��O_*_2S  !8_@[L �O�_C#�O �_
_�_�_@_�_d_v_ ?o�_Zo�_jo�ooo o*oDoNo�oroD V�oz�o�o|& ��
�n���� :��������"�ʏF� X�!�|�<���`�r�֏ ����L�՟0��T� � &�8���D���ҟ�^� ���گ�P��t��� ���4�ί������� (�:��^�ς�B�T� ��j�ܿ����6� ��ߎ�~ϐϢϼ��� @��ϖ߼���2���V� h�z��ߞ�J�p���� ��
��.�� �d�$� 6���B��������� �����N� r���M ��h��x��� 8J\��,Rd ������F //|$/��{/� �/��/�/0/�/T/f/�/?�4S�2�?4:ψ  �B4: 8�1�?�)
 �?�?��?�?c:UD1:�\�<��F1R_G�RP 1�K?� 	 @� :O LK6OlOZO�O~O�O�N��@�O�J�A�?_�O<7_"U?�  R_d[ N_�_r_�_�_�_�_�_ �_�_&ooJo8ono\o0�o�o�o�o	5�o��oD3SCB 2P; =_:L^�p�����:<U�TORIAL �P;�?�?7V_C�ONFIG  �P=�1�?�?t�$�OUTPUT !P9e�����ď֏ �����0�B�T�f� x�����b���ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϷ� ������ ��$�6�H� Z�l�~ߐߢ߳����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� �����&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/N�`��� �/??&?8?J?\?n? �?�?�?�?�?��?�? O"O4OFOXOjO|O�O �O�O�O�?�O�O__ 0_B_T_f_x_�_�_�_ �_�_�O�_oo,o>o Poboto�o�o�o�o�o �_�o(:L^ p������o�  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�nπ�ϒϤ϶����Ͻ(���������� 6��/Z�l�~ߐߢߴ� ��������� �2�� V�h�z�������� ����
��.�@�Q�d� v��������������� *<M�`r� ������ &8I\n��� �����/"/4/ F/Wj/|/�/�/�/�/ �/�/�/??0?B?S/ f?x?�?�?�?�?�?�? �?OO,O>OO?bOtO �O�O�O�O�O�O�O_ _(_:_L_]Op_�_�_ �_�_�_�_�_ oo$o 6oHoY_lo~o�o�o�o �o�o�o�o 2D�S{�$TX_SCREEN 1"�����}�S�������Bք1�C�U�g� y�������ӏ��� 	����?���c�u��� ������4��X��� )�;�M�_�֟蟕��� ��˯ݯ�f����7� I�[�m�������,� ٿ����!�3Ϫ��� i�{ύϟϱ���:��� ^���/�A�S�e�������$UALRM_MSG ?sy��p ��Vj���� ����"��F�9�K�i�o���������S�EV  ������ECFG �$su}q  �Ve@�  AJ� �  B�Vd
  ��]csu}��������� ������1?&�GRP 2%0�; 0Vf	 g�����I_BBL_N�OTE &0�T��l]b�xp_a<�DEF�PRO��Z�� (%��_`�* N9r]�������/�FKE�YDATA 1'<sys p ?�Vfvy/�/b/�/�/�*�,(�/�/Vd([ INST ]�/��.  IRECTR�D?+?ND=2T?V? CHOICE?��?[EDCMD��?�?� ORE0FO�?�?O*OONO5O rO�OkO�O�O�O�O�O�_�O&_8_ ���/frh/gu�i/whitehome.png9_`w_�_�_�_�_�PVinstb_�_oo�(o:o�W  QUdirec�U�_o�o�o�o�oVhinaj�o�);�oXfchoicaS�o�������PPVedcmdo��'�9�K��V}PVarwrg�o ��������ϏVx��� �"�4�F�X��|��� ����ğ֟e����� 0�B�T��x������� ��ү�s���,�>� P�b�񯆿������ο �o���(�:�L�^� p�GUuϜϮ������� �����,�>�P�b�t� ߘߪ߼������߁� �(�:�L�^�p��� ��������� ���$� 6�H�Z�l�~������ ����������2D Vhz���� ��
�@Rd v��)���� //�</N/`/r/�/ �/%/�/�/�/�/?? &?�/J?\?n?�?�?�?�?[�;�JP����?�?�=�? O2OF,_cO_�OnO �O�O�O�O�O__�O ;_"___q_X_�_|_�_ �_�_�_�_o�_7oIo 0omoTo�o�o���o�o �o�o!0?EWi {���@��� ��/��S�e�w��� ����<�я����� +�=�̏a�s������� ��J�ߟ���'�9� ȟ]�o���������ɯ X�����#�5�G�֯ k�}�������ſT�� ����1�C�U��y� �ϝϯ�����b���	� �-�?�Q���u߇ߙ� �߽����߸o��)� ;�M�_�f߃���� ������~��%�7�I� [�m������������ ��z�!3EWi {
������ �/ASew ������/� +/=/O/a/s/�//�/ �/�/�/�/?�/'?9? K?]?o?�?�?"?�?�? �?�?�?O�?5OGOYO kO}O�OO�O�O�O�O��O__��![�>�����J_\_ n]F_�_�_|V,�o�_ �o�_�_o-ooQo8o uo�ono�o�o�o�o�o �o);"_F� j������� ��7�I�[�m�����O ��Ǐُ����!��� E�W�i�{�����.�ß ՟�������A�S� e�w�������<�ѯ� ����+���O�a�s� ������8�Ϳ߿�� �'�9�ȿ]�oρϓ� �Ϸ�F��������#� 5���Y�k�}ߏߡ߳� ��T�������1�C� ��g�y������P� ����	��-�?�Q�(� u��������������� );M_��� �����l %7I[��� ����z/!/3/ E/W/i/��/�/�/�/ �/�/v/??/?A?S? e?w??�?�?�?�?�? �?�?O+O=OOOaOsO O�O�O�O�O�O�O_ �O'_9_K_]_o_�__ �_�_�_�_�_�_�_#o�5oGoYoko}o�of���k�f�����o�o�m�o �f,�C�gN�� �������� ?�Q�8�u�\������� Ϗ���ڏ�)��M� 4�q���b�����˟ݟ ��o%�7�I�[�m� ��� ���ǯٯ��� ���3�E�W�i�{��� ���ÿտ����� ��A�S�e�wωϛ�*� ���������ߨ�=� O�a�s߅ߗߩ�8��� ������'��K�]� o����4������� ���#�5���Y�k�}� ������B������� 1��Ugy�� ������	- ?Fcu���� �^�//)/;/M/ �q/�/�/�/�/�/Z/ �/??%?7?I?[?�/ ?�?�?�?�?�?h?�? O!O3OEOWO�?{O�O �O�O�O�O�OvO__ /_A_S_e_�O�_�_�_ �_�_�_r_oo+o=o Ooaosoo�o�o�o�o �o�o�o'9K] o�o��������� ��� ���*�<�N�&�p���\�,n���f�׏ ������1��U�g� N���r��������̟ 	���?�&�c�J��� ������������ )�;�M�_�q������ ��˿ݿ�ϐ�%�7� I�[�m��ϣϵ��� �����ό�!�3�E�W� i�{ߍ�߱������� ����/�A�S�e�w� ������������ ���=�O�a�s����� &����������� 9K]o���4 ����#�G Yk}��0�� ��//1/�U/g/ y/�/�/�/��/�/�/ 	??-???�/c?u?�? �?�?�?L?�?�?OO )O;O�?_OqO�O�O�O �O�OZO�O__%_7_ I_�Om__�_�_�_�_ V_�_�_o!o3oEoWo �_{o�o�o�o�o�odo �o/AS�ow ������r� �+�=�O�a������ ����͏ߏn���'��9�K�]�o�F q�}�F �����@���������̖,ޯ #�֯G�.�k�}�d��� ��ůׯ������1� �U�<�y���r����� ӿ����	��-��Q� c�B/�ϙϫϽ����� ����)�;�M�_�q�  ߕߧ߹�������~� �%�7�I�[�m��ߑ� ������������!� 3�E�W�i�{�
����� ����������/A Sew���� ���+=Oa s������ //�9/K/]/o/�/ �/"/�/�/�/�/�/? �/5?G?Y?k?}?�?�? x��?�?�?�?OO&? COUOgOyO�O�O�O>O �O�O�O	__-_�OQ_ c_u_�_�_�_:_�_�_ �_oo)o;o�__oqo �o�o�o�oHo�o�o %7�o[m� ���V���!� 3�E��i�{������� ÏR������/�A� S��w���������џ `�����+�=�O�ޟ s���������ͯ߯�0����0���
��.��P�b�<�,Nϓ�FϷ���ۿ �Կ���5�G�.�k� RϏϡψ��Ϭ����� ����C�*�g�y�`� �߄����߲?��	�� -�?�Q�`�u���� ������p���)�;� M�_������������ ��l�%7I[ m�������� z!3EWi� �������� ///A/S/e/w//�/ �/�/�/�/�/�/?+? =?O?a?s?�??�?�? �?�?�?O�?'O9OKO ]OoO�OO�O�O�O�O �O�O_��5_G_Y_k_ }_�_�O�_�_�_�_�_ oo�_CoUogoyo�o �o,o�o�o�o�o	 �o?Qcu��� :�����)�� M�_�q�������6�ˏ ݏ���%�7�Ə[� m��������D�ٟ� ���!�3�W�i�{� ������ïR����� �/�A�Яe�w����� ����N������+�h=�O�&PQ��&P���zόϞ�v����Ϭ�,��߶� '��K�]�D߁�hߥ� �ߞ����������5� �Y�k�R��v��� ���������1�C�"_ g�y���������п�� ��	-?Q��u �����^� );M�q�� ����l//%/ 7/I/[/�/�/�/�/ �/�/h/�/?!?3?E? W?i?�/�?�?�?�?�? �?v?OO/OAOSOeO �?�O�O�O�O�O�O�O �O_+_=_O_a_s__ �_�_�_�_�_�_�_o 'o9oKo]ooo�oX��o �o�o�o�o�oo#5 GYk}��� �����1�C�U� g�y��������ӏ� ��	����?�Q�c�u� ����(���ϟ��� ���;�M�_�q����� ��6�˯ݯ���%� ��I�[�m������2� ǿٿ����!�3�¿ W�i�{ύϟϱ�@��� ������/߾�S�e�@w߉ߛ߭߿ߖ`�����`�����������0�B��, .�s�&���~����� �����'��K�2�o� ��h������������� ��#
GY@}d ���o��� 1@�Ugy��� �P��	//-/?/ �c/u/�/�/�/�/L/ �/�/??)?;?M?�/ q?�?�?�?�?�?Z?�? OO%O7OIO�?mOO �O�O�O�O�OhO�O_ !_3_E_W_�O{_�_�_ �_�_�_d_�_oo/o AoSoeo�_�o�o�o�o �o�oro+=O a�o������ ���'�9�K�]�o� v������ɏۏ��� ��#�5�G�Y�k�}�� ����şן������ 1�C�U�g�y������ ��ӯ���	���-�?� Q�c�u��������Ͽ ���Ϧ�;�M�_� qσϕ�$Ϲ������� �ߢ�7�I�[�m�� �ߣ�2���������� !��E�W�i�{��� .�����������/���$UI_INU�SER  ����P���  0�4�_M�ENHIST 1�(P�  �( ]����(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1o������)����631��ew��� �'-?7@S��
��.��?edit��SO�LDADORA,A3!t����35�GMAIN_XU@_��/ /��,��GIR_HOME �x/�/�/����/�/ �/�/??,?�/P?b? t?�?�?�?���D1�� D?�?�?OO)O;O>? _OqO�O�O�O�OHO�O �O__%_7_�O�Om_ _�_�_�_�_V_�_�_ o!o3oEo�_io{o�o �o�o�oRodo�o /AS�ow��� ���?�?��+�=� O�a�d��������͏ ߏn���'�9�K�]� o���������ɟ۟� |��#�5�G�Y�k��� ������ůׯ����� �1�C�U�g�y���� ����ӿ�����-� ?�Q�c�uχϊ��Ͻ� ������ߔ�)�;�M� _�q߃ߕ�$߹����� �����7�I�[�m� �� ���������� �!���E�W�i�{��� ��.��������� ��Sew��� �����+� �as����J ��//'/9/�]/ o/�/�/�/�/F/X/�/ �/?#?5?G?�/k?}? �?�?�?�?T?�?�?O�O1OCO.��$U�I_PANEDA�TA 1*����yA  �	�}  fr�h/gui�Ade�v0.stm ?�_width=0�&_height�=10�@�@ice�=TP&_lin�es=15&_c�olumns=4��@font=24�&_page=w�hole�@UO1)�  rim�O!_  �@8_J_\_n_�_�_ �O�_�_�_�_�_o"o 	oFo-ojo|oco�o�o��o�o�o�o1� ��     I}�2_7I [m��o�(_� ���!�3��W�i� P���t���Ï���Ώ ���A�(�e�w�^���y��{C�۟� ���#�5���Y��}� ������ůׯ>���� ��1��U�g�N���r� ����ӿ�̿	��-� ?ϲ�ğuχϙϫϽ� ��"���f��)�;�M� _�q߃��ϧߎ��߲� �����%��I�[�B� �f������L�^� �!�3�E�W�i���� ����������� ��A(ew^�� �����+ O6s������� ��//h9/��]/ o/�/�/�/�//�/�/ �/?�/5?G?.?k?R? �?v?�?�?�?�?�?O O��UOgOyO�O�O �OO�OF/�O	__-_ ?_Q_c_�O�_n_�_�_ �_�_�_o�_)o;o"o _oFo�o�o|o�o,O>O �o%7I�om �O������ d!��E�W�>�{�b� ������Տ������`/��S��o�o}�d�@������ӟ���)�� ��u�H�Z�l�~��� ��	�Ư���ѯ� � �D�+�h�z�a������¿Կ�����x�c�k��$UI_POST�YPE  �e�� 	 ��[�*�QUICK�MEN  9��H�^�,�RESTO�RE 1+�e�  ��뿑r�����ϑrm  �)�;�M�_�q�ߕ� �߹����߀���%� 7�I���V�h�z��ߵ� ���������!�3�E� W�i�{���������� ��������Se w��>���� �+=Oas (����// '/9/�]/o/�/�/�/ H/�/�/�/�/?�? 0?B?�/}?�?�?�?�? h?�?�?OO1OCO�?�gOyO�O�O�Oi�SC�REy�?~��u1sc��uU2�D3�D4�D5�D�6�D7�D8�A�CT;AT5�� ���e"�USER�@�O�B�T�@�Cks�C�T4��T5�T6�T7�T8��Q*�NDO_CFG ,9�t�s�*��PD-QgY�None *��^P_INFO 1�-�e`��0% �O,o�xo[o>oo�o to�o�o�o�o�o!�EW:{b��QO�FFSET 09�a�PC��XO� ���/�&�8�e�\� n��r�����ȏ��� ��+�"�4�F����ϒ�Ā���
��ڟ�xUFRAME  PD��V�QRTOL_�ABRT���s�E�NB��GRP �11�Ɋ�Cz  A�u�s��Qs��� ������ͯ߯��x��U?��Q.�MSK � B�a.�N���%	i�%b���k�V�CMR[�27�{S#�R@	�Pfr�1: SC13?0EF2 *ݿ��PD�����T&��5ZR@�Q?��@�up��ȇ� ɟ5�?�IH`�rϟ�ıh����8��A�RB����RB B����RA#ի�D� ��h�7ߌ�w߰ߛ��� ����
�a���@�+�=��v�)ߚ�ISI?ONTMOU�B���U���R8�SﳸS� �j� FR:\���\�PA\�� ��� MC�L�OG�   U�D1�EX5�RA'� B@ ��x�I�r���I�����PC � n?6  ���IFu��%��`��Z�  =���PD	 �J�*�TRAINp_���ǐ  dP�p	�栲9�}( c��W���� ���.2@R�dv���_\�RE���:b�ʲ��LEX�E��;�{�Q1-e~��VMPHAS/P��U�SЖ�RT�D_FILTERw 2<�{ Ԓ��,�{/�/�/�/�/�/ �/�/??��i/N?`? r?�?�?�?�?�?�?�?���SHIFT�1==�{
 <��q� JODU)OOO�O_OqO�O �O�O�O�O�O_<__�%_r_I_[_�__	�LIVE/SNA�Pesvsfli�v.�_��� �pU�P�Rmenu �_�_�_Woio@b	E��>IO�EMO��?��� ��$WAITDINEND��+��dO?�"��g���o�S�iTIM@���<|G�o^}�o�{�az/azN�hRELE%!@��d�����a_ACT�P�K�E�� @d�ko���E�RDIS�PA��`�V_AXSR�p2�Ab�����Vp_�IR  �j  	��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i�{�������ÿ�տ�������XV�R�aB��$Z�ABCp1C�� ,N f�2ϵ�Z[IP��D�e�������ύ�MPCF__G 1Eٍ0J��=��S�FىX�`#� �c�߆�<90 �߻�S�|��ߠ�?�}������ S��$�z�8���� ���������@��
�4�M���G��|JÛ�YLINDK!�Hً Є� ,(  *������`���������� �� );M��p���{ ��� U6 ��lS�w������Y�2Iه]� �)�#/3,���\/@G/�/��/�/���!�A�c�SPHER/E 2Ju��*? z�/<?#?`?��/�? �?$�?k?Q?O�?&O O?\OnO�?�?�OO �O�O�O�OEO"_4_F_6M�ZZ/� ǘf