��   F��A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A #  �����#�AMON_D�O_T   �$PORT_�TYPE  �@NUMJ/SG�NL7 L�$MIN_RAN}GI$MAXr�NOo ALxp V��~ �COUNT>J �AWE08 �� $AWn0ENBJ $�|G1LY_TIV�$WRN_ALM�STP�
�E��C�.�WT�C�
J�AFT_�CHGxAVRG�_INT��{SgAVE�YP1?ER_REG�Tw$WA� SIG�� OP��V/OLTS�����AMP�&AEx �#E_VL� �&D'>% I*f$� _�ANL�  �p 
$US0 S�_CMD � PRIORITY�"�UPPER� $�LOW�$�#$FgDBK�"�RAv ~�!SQ_AVG�#n�#SD_� CE� r� ��$ �� � LIN�!$A�RC_ENABL��!� 0DETEC��!< ELD_SP~�$PD_UNI���!92DIS�"�I�D IM�#���  v1WFt2S_�P�CF�" �� $PS_MANUF �2�ODEL�5PRO�CESN0�0WFE�EW0ESC�2�2_�FI#1�1�1�7T _SAO�"�2I�6D�7�DC1�6L �"{2 �� CNV� 7   $EQ��zxODOU���?@TBd� �$?C 2 �Y>ADD   �, � MM�!�$D� ��!?2 $F� �B�?@7	JBSEL�10_NOJDAT�A_s@�@  V�WPpG
{M
{"v�AWP7 L@��L
 �WIR�_CLP4 �L@ASBU8  HG $4���R�4�YPREFx� �U�1_ECU���  JB~ �S �  $BPEtEPf#}!SCH7 � �!��``�1e#dPK*j�FREQ.gULSwbSP�0fg2y��!hyb*g�F�AI6 �ZCoVG }�hp dD�e�e�`�	��a��dBVB�aZ�EROy}uSLYO]R�`NT�!P�c�O	U\93�L FORMA0NAra�0J3W	� D�cQW�UXWEIOEX>74 �A�iWfxccpS_91INp� :1�U�p�� FAUG"t0LIO�0�qP�!�G���R<�ADp;�STI�C�@�pROBOT�ADY�rERRMO�SE��`S���p�!TR��$S�CHDOG_�@%��0?_ACTIV���UI�C�01�2�q�OTF7 � $
��P��x0�nfpNCi0� c;�f0�*d;�*g0� 7f;�7i0�Fd;�Fg~�Td��TfUP�@�B?P� PCR7�� WSTK��� =�Hr ՒƁ%��00���2�X���0A~�3KIPTHE91�S;�8�����PIKEf��p�0�0WWV�2t�E_HO;0�0���PHK-1���� R�MT���SPTL��0p�$Hz��SyW��pd$BBg1�_ONL4�$B��2pf�bgF�WF �1e2_R��zE"�!� �_W;6�AND1OsFF���!ND2g�	3g�R�S� �A� �t�PM� | $�0�@g��e��*f���7b��Ff�TfAD�APT� G�CSENS�c��!ݒ��8 � 0?,2�� �"��$�1b�!c�7c c�Fa|�Tac�^��'y�P�&l��&�!4�&5�&�6�"8�W�@�2 HOEU�!�o � �SE�0�g4�Q�T <��6�'��46�q56��0� %$CUR�R7(��"HEATzPe@�!燰"j����i�p��GAP�#Ti�XPY0��EHP��@�f�pDS�@�!GP�0�S�!$���$GOf� RI���AM�#$/"�#M��jAN3O�'BEFB ;�LHV1 [5j��43;1 `H�V�!PA�H�r���3��F10�� �c2�SR 7_ � 	� RSB�$��0G�m�b�O�J���O��DU�IDW�AXQl�2C,1�L�"D����?3��R9G�8  4�@P��q]ִSGʦ�~�;A�8�8  $ $��@�CL�$��s	�<y��$ ; o2� �"�ql��q��� 	PK�P��
��* ���q�Ba��b*�@4�5�6:2�K�3�����FW��q�B��ALAR���2��2������
�3�Q_R }��
�.44�F�+�PW,���_@ĸ�� �]�������Q`bwm��t���QDI��c�j��~pus�R�S�IZ���BOAR����1]E7�]�@\�h"0h"��ľ��$VEND��I>��DEVIC��0�D����MAJ��V�#IN�(�$�uI"�vcMA��pFI�0�BW�ۓ�� p $��X�� ⡡��MF̀OR_R��C��^1D4TO_��O5_�R�pRS�Q'�OS�9�rUP� #N��S�0�`�=� �6��6��9PUR�G��RKtSTFR�p&���A��.E��.E�AED��P-��M�%�fMT�����eEM 7��Q�5���Z$�22��9�P駇��K�p�QAsDJ�T��NEXT�N�r_LE�c��P��X��M����aA��!_�#IV���H�q�2F�eFL������P�†U���0�8� ��TW�T[�CY�� |���  �	`�`( �bTOTACL_�Q�c���VI�p��WWARo��U��A�*�PY&1b�uK�G���'" A}�#Nޓp  �aSC�FG�1z�LCOO�B:��P�Q��S!@���GLOB��P�⣠� ��NOT��$0QI4�*��AVh�Y��$���������e��W_SH�FL�W�X�fkrI`�$�q �e�RY	���оP��%�ʀLIM�S`�i�@�c7�UIF��e�APCOUP}L�R @ �pؓq��� �qUR�`N��<�MMY`m �u0�u�  ��ޏ�USTOk�    x�0 �q�p` 
!3SEM�Gg��1! ,��M�G�Ag���NOzPR� ����wa�"� ,/���Ȣ=6Ƞ��3T� )�RT���p�`��=����AHER� ��A�������'"݈{ �������@���Q�L� �)BD ��2C���7B�<�i3_FIL@�Wn��BUG_3SM ���ñF_F����q�4, _4N SV@БT�C�P��=Ҕ�DIO�������.a�3TM�C��PA�Pq���qw�x��q�_DY�NV�2Wԣ����KEYV�GQׂ���F��?�/B�{�_C:��R�TOU����8�Б��CAL�Q0D�`� TIp1�P_y��RT���@��A?2��$$CLAS�S  ������ ��� �-�S�B���  ����IRTUx�����AWAOY1��� 
��$�a
�K���n�2�f�[�[���g�
�?�������g��� ��������(�:��L�^�pςϑ�l�EXEu�`���������Ͽ �*�<�N�`�r߄ߖ�p�ߺߕ�r@S Rw���:����#�5�G� Y�k�}���������������l�NLG7 2x� �����E?��<1�6�`��e�� p`����{` 2�:�)��General Purpose��MIG (V�olts, 0)���� ����
AW�MGENL.VR�A*EGLM#G19��g�`�� ������'���������������C�NV 2	x��[����� 4aPzUh �����//� =/O/./s/�/\�/�/ b/�/�/�/?'??K? ]?<?�?�?r?�?��E �/�?O�?2ODO#OhO zOYO�O�O�O�O�O�O 
__�?@_R_�Ov_�_ g_�_�_�_�_�_�_o �_(oNo�?ro-_�o�o 3o�o�o�o�o8 J)nM_�{o� ����� �F�%� j�|�[�������֏� go���0�B�!�f�E� W���{���ҟ����� �,�>��b�t���� ����ί௿����� :�L�+�p����O��� ʿU�� �߿$�6�� Z�l�KϐϢρ����� ����ߵ�2�D�#�h� z�Yߞ�}ߏ��߳����
��NVWP 2�|	i\>�T 
���b�t���UST�OM 2|l  ��������h��	hd"���DEF�SCH R|��Q�<�b�@De�fault Schg���n��������� ��K"4� Xj��������
)�FBKLOG�1 @��T���  Ugy��12=O�����5LG_CNT � ����)�IOE�X 2�����A� ��C�]$@�������!�
Weld Spee%�~�IPM  d$ �/�/�/�/??(?:?~��OTF 2���A?�?�?�?�?�?�C8=�����@����?K)�PCR k2��pI�BH�?��BC!�FK<D7�������?�ffA�Z �A"��OFM"@�����/�O@O�"@�����WOELG��k%*_�F��0234567O8901JRUK%4_y_�_�_HIȩ_7]�O_OSRAM2��I�B�$�_oCRGS_EL R<�Q�� 	Proce�ss 1oSf2T�_oj3i�o4i��o5�-mlXS��R�o7��kn8i'l�"@��� �_);Es-B� �W�%�Volta+ge��qsfc%�Dw|!@]y��h��aWiore f�  s�$	� hc%[&t/�o DS�l*�<�N�`�r� ��������̏ޏ��� �&�]+zvd"�����  �#��E��Z"!��a��^/�� ��V���a�aɒ�Curren=t�Amp�=� ��l�eu���Q�c�u� ��������ϯ��� �)�;�M��W���a�� ���ឱ	q��)q��Iq ��R�͹ϧg�a�aA� �b-���-�	q-�)q-��VE!��\e�	q/?�����Z�%�� ����ϻ������PD�RuS R\zH�� jq��C�U�g����� gߩ߻�u߇ߙ��� ������]�o�)�;�M� ��������#��� ���k�}�7�I�[��� ��������1C�� I��Wi�� ����?Q /������/ /)/;/M+�U/g){/��/�/M/�/?cS2�S�^=R��b�S2UP�Yp^=�=�o�?�33H1>E0=OL��>I0h!�"�#�$�1t9�g��q�#?�v�#>��8�8CWIRE �2&M<�?�?h��>�3�>�G(�=�J*�ESCFG �G�A��Y���OOˎE7])COU�PL�0=k
0 �vkB`�D�^�L�[�O ZW�O�G_�OP_G_Y\>�HNB  ��Ec�&FUSTOM � =k
8ƙy�O&EE�MGOFF !�=kS��)BPCRg "�_�@���zqC{sUūMJo�\zt�f_oeo��
Cl�q� �1