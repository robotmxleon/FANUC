��  X>�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A3  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ���AIO_CNV�w l� RAC��LO�MOD_T�YP@FIR�H�AL�>#IN_O�U�FAC� gINTERCEPf�BI�IZ@!LRM_RECO"w  � ALM�"�ENB���&ONܢ!� MDG/ �0 $DEBUCG1A�"d�$3A�O� ."��!_IF�� P $E/NABL@C#� �P dC#U5K�!M�A�B �"�
� O�G�f d PC�OUPLE,  w $�!PP_D0OCES0�!e81�!�f R1> Q� � $SOFT��T_IDq2TOT�AL_EQ� $̋0�0NO�2U SP?I_INDE]�5�Xq2SCREENo_NAM� e2/SIGN�0e?w;��0PK_FI0	$THKY#GoPANE�4 � �DUMMY1d�JD�!UE4RAG_��ARG1R� � $TIT1 d ��� �Dd�D� �DTi@�D5�F6�F7�F8�F9�G0�G�GPA �E�GhA�E�G1�G ԈF�G1�G2�BME��ASBN_CF��!	 8� !J� ; 
2L A_CM�NT�$FLAsGS]�CHE"�� � ELLSET�UP 
� $�HOME_ PR�<0%�SMACR=O�RREPR�XD0D+�0��R{�T �UTOB U��0 9DE7VIC�CTI�0�A� �013�`B�S�e#VAL�#ISP�_UNI�U`_D�ODf7{iFR_F �0K%D13��1c��C_WAqda�jO�FF_U0N�DEL�hLF0EaA�a7b�??a�`$C?���PA#E�C#sAT�B�d��0W_PLv�0CH/ <� PU�P�B
2ds�`�QgdsDUT�P�HAgpSF���WELDH2/�0 =Lc7w7atAING�0$�r�1�@�D2�4%$AS_LKIN;tE�w�t_�~�2UCC_AS
B�FAIL�DSB�"�FAL0�AB<�0�NRDY��P�z$�YN�Wq<��`DE6r��`���p+�����tSTK��0+�;s7�;sNO�p��[�̈́r��U* Ȁ%� 9 � �� ��q`�G�pC�G�+�U�S_FT�0vpF�ǂG�SSF���PAUS���ON\7xǓHOU�ŕ�MI�0�0ƔSECȲ2�ryi �rHE8K0�v8vGAP�+�r	�I� � GTH�F��D_I���T=  �l�����`�s9!̅0����9!G�UN1����q���#MO� �cE' � [M�c�\���REV�B7�~����AXI� ~�R  � sOD�P-��dPM�^Q%�;�/�"8�� F�q��!X�0DfT p{ E RD_E%�~Iq$FSSB�&_$CHKB�pEde#AG� �p�  "
�$Ա� Vt:5���3�
`a_EDu �� � C2��qS��`�vl �d$OP��0�2�a<�_OK<��Y�TP_C� <�pd�vU �PLAC��^}��p� xaCOM	M� �rD|ƒ��0�`��KO]BMpBIGA�LLOW� (tK�w�0VAR��xd!�1�q�BL�0S � ,K|a�r�PS�`�0M_O]|=՗�CCG�`=N�! �� ��_I_��� �0�� �B.��1S� ~�CC'BDD�!��I����0�@��84_ CCWp` OOL
��P'�M�M
�n�CHs$MEAdP�d`T�P�!���TRQ�a�CN���FS3��ir�!/0_F��( D�!��v CFfT X0�GRV0��MCqNGFLI���0UJ�p����!� SWIl��&"D�N�P�d��pM~� � �0EED��!��wPo��`�PJedV
�&$�p��1``�P��ELBOF� �=��=�p/0���3P�� ���E���G� �>A0WARNM�`ju���wP��𼠤 CO�R-�8`FLTR^juTRAT Tlp�� $ACC�rT�B� ��r$OR1I�.&��RT�P�p�gU�HG@I��"3�T{�1�I �rp������ ���0�"�Q���HD���a
�2
BJ{PC��U3�4�5�6��7�8�9��COfS_rt����3�V�OLLE�C��"MULTI�b
2��A
1;�0�T_�R  4�� STY2�R���).��p�b�n� |A06Kb�Ib�$���Pc���UT�O=�cE�EXT�!Y�
B!�Q O2 
l��a0��Ru�r����  �"���Q�@���qc0n~#!|��1Y�M
�P8$�  lTR�� " Lq��/��P��`AX$JOB`׍���4IGx# d��?%?78���3�p%��u�� _wMOR��$ t���FN�
CNG&AF�TBA���6�JC���9��D@r��1CUR�.KPa`/E;��%��?��ttaoA��XbMJ��_R��|rC�LQJ�r�H�LJ�DA����I�����2G���jRfT&� ���bG���HwANC6$LG�� iqda��N�*�YaCᇁ��0|rf�R'L��0mTX���nSDBWnS3RA�SnSAZ�P�Xp��$  ' FCT�іe�_F��Pn�e�M
P�QIkOh��� ���1��e���Cg�0��A���MPa� 6��HK�&AEUp�p��Q�A 9 �' � ]PI��CSsXC��Zq( xs���s��T�R�CcPN콰��MG�IGH�"��aWIDR�$cVT�P��9�EF�iPA cI�XP,a|Q�1u�CUST��uU��)R"TIT�4���%nAIO��x �BG_�L���*c \q���OR��@$!�q���-��OeP ��jЅpIp�Q�u�J�8�
��0��DBP_XWORK��+��$SK0����1D�BT)PTRw� , �l@Ab��s�R�0�ؠD��A:0_C`����=�+`H�PL�qD��R�A�"��#�D���r�����BJ���9l��� X@DB�Q2��-�r~qPR��ΰ�
�ct��. p�E�S�a�
�LӉ�/��b���( ��0��b��Pj� 91%�7�ENE��0� 2D�7���RE\���3HPC� � .$L��/�$Ӄ�����INE�׶�q_D����ROS��E0"2q��f0��p��PAZ�tAsbE�TURN����MR�Q2UA@�CRŐE�WMwp��SIGN�A&rlPA��W�`�0$Pf13$P�P�2j���!q������DQ���f������׶GO_AW;0���vp��qa��pCS'���CYx42O�1�8�8�*��2��2�N�@�x�CtDۣDEVIѐ� 5 P $�RBֳ��I�P<.�i�I_BY�q��T�A9�HNDG�6�������b�DSBLr3ͳ��ςݡLe7 H� �� ��TOFB̶�FEБg')�h�ۣ�f8��DO�a�� MC9�"�`�s(r�(��H�PWp���ܢSLA4���9IINP!Ѐ� ж�|ۡ�:D *�SPNp�#�lƍ�1��W�I1��J��Eȅq87�qW��NT�V#��V ��SKI�STE^��b��p�L��aJ_�Sjb_>����SAF�k���_�SVBEXCLUT��po�D�pLX ���YH��%q��I_yV9`�bPPLYj���������_ML���L�VRFY_4D��M�IO�`   P�%`�b�Oe��LS�|b��4}�$�����P�u��l�Y�AU NFzf@�����)���cD�4dͰ� S��r�AF� �CPX���&`� 3;j��pTA#����  
�i�SGN��<��<@3�P��c _�t�a���qd��rt��`UN>�����<@rD�p]�T`����%`X����zrEF�pI>�= @��F��\t6@OTS����|�����h�塁x!Mr�NIC!>2K�GM A��i�DAY�sLOADЩ��D��5�� �[EF pXI�?j����~cO� �5�_�RTRQU�@ D�����0Q�p B�EԠ��� ?K�%>`� ��AMP*Pp��A�"'; DB�'��VDUS�U�.�CABU�B`��NS9@ID�1W�R$�Q!`V[�Vq_#� ; �DI@�J$C� /$VS�SE�T�BDC�A�� ���|�DB�AE_l�;VE�P�0SW!�!�@x�3�2� @�`�OH�@3PP <IRwqDBB�p�=�!U����t"BAS��o'~P�Pn%[�d� B	� ����RQDW]%MS�� �%AXC'�;LIFEC���� ��	2�N14B5��34BChd@/Ź�Cq`ʡaN�4q�6��OVՐ�%6HEh�DBSUP$�1��	2D�_�4j�BH1_!C�5š�7Z�:W�:qa�7�S��"BcXZ�Pʁ4AY2HEC��T�pސ�NM���
�0P�dD `�L��@HE�VXCSI�Z?6k0��[�Nh�U7FFI�0��C���������6����M�SWJEE 8��K�EYIMAG�TM���S�A5��F��
q��Y�VIE �qF 	�PLQ�_�ӛ?�@A�D&`KDG�� ��ST��! >R|�FT��FT� FT� >FPEMAILb �xaA���FAULS�HR�*�;pCOU�_��q�T��U�IO< $�S_�S#v�ITճBUFkG��kG@�jp`p�0B�Tk�C��Rws�PSAV(e�R�+Bd�$ Cg�p��P/d_ň��$̰_�Pec �iOT����P@����jA�gAX�sq:p�P���\c_G3
I YSN_e!�pJ0Df�TW�r�d"MO_0T��F��� 2���$^ЈqK��ey&^��5r�)�4��qL�0��nq�S�cC_ܐ��AK씐pu�t��R�A8�u�XnqDSP�FnrPC�{IM5c�s�q�nq�U�w{0�0�F�PIPR�nsN!Djp��sTH��"ûr� T�ߑ�sHSDI�vAGBSC_�9@`�V���x�v��c~����NV���G��~�*@�v�PF�!�`d�s0p�a��SqC�\��sMER��>nqFBCMP��mp�ET�⌐M�BFU�0DU�P?�M�B
�CD�yH��`�S� R�_NO�ዑN� `%�i�cg��PSf��Cjpv�C���ap*Qd��`U OH�� ��c d�������}� 锍��9疗疢�疮A�7�8�9P�0��1��1
�U1�1$�11�1>�U1K�1X�2f�2���2
�2�2$�2�1�2>�2K�2X�3Jf�3�3��
�3�U3$�31�3>�3K��3X�4f�~QEXT�TP <sK�p@<6p�p2ǋ��`�FDR�QT�PV��b	2p�v�	2�REM�F��0BO�VM�s��A��TR�OV��DT3`��MX��IN��Q0�ʶ'IND���
	�i��`$DG�a{#���4P5�D���RI�V"�=20BGEAR��qIO�K��;N 0p}ة�(���@�0<�Z_MCM@	1_��F|0UR"�R y,t� a? P0��?��!?��EG��jqa��e©S� � P�a�R�IM���SETUP?2_ T � �STD6���<����I��C��Ո CrU T([ �RTt)Nz%��+p�IFIQ!+p���А��PT{b*QF�LUI1TV �3 Y�PUR�!遀W2�r<qv��P�� I��$�S��?x�#�JQpCOw`�cV�RT� x$SHqO���SASSY���a?58������AZ�W�RFU��15q:��25qine��*@�X |�NAV�`��3���*@x�R=1��VISIJ�&��SC���E�c�T\�AV��O���B%EX$P�O��I\ ��FMR2b�Y o�X�}p�bpN t�{ߍߟ߶ơP���%_f�G�_��B���M4�Y�k�DGC{LFR%DGDYLD��7�5!6.�04R��MR�3SZ�@�	? T�FS�`2T�[ P!��bs�`�$EX_���1P�`Ā\2�3�5�S�G��9\��
����PWeO�&DEBcUG��"��GRR�spU�BKU�O�1�� 0PO@� ;)' ��' Mb�gLOO�ci!SM� �E7bjq��� _E �] �@Y�*QT�ERM�%^�%v�O�RIBq� _�%��S#M_OpL� `�%1d���(a�&��UPR�b� -���Q]�#0^��G:�0ELTO{Q$wUSE��NFIc1�G2��!���$4_�$UFR��$`j�A1}0=�� OT�7ƭ�TAX�p��3NSTCpPATM�d@�2OPTHJ�;�E4P8_bD�H2ARTP`R5p�PPa{RG1REL�:�aSHFT?�H1�1��8_N�R�8��& � $�'H@a�q�B���bSHI@�Uz�� JaAYLO� �a�a���Y�1��~�J�ERVA�3H 7Cp�2�����E����RC�~�ASY1M.q~�H1WJ[7���E��1Y�>�U�2TCp�a�5�Q=��5P���@��bFORCpMLKa�GRz!:c���'"`&�0w0�a�HOb�fd Ԟ2��& �X�OCA1E!��$OP����V�t F����P��P��2`RŃ�aOUx��3e��R�5Ie h�1���e$PWRL�IM;e�BR_�S�4��� �3H1UD�kp�Q�Bte7�$HSu!^�`ADDR2�H}!AG�2�a�a�ab�R��.x�f H!�S��񀌳u��u
�u�SaEv��Y�w�HSH�;MN��g
 �P0r��T�@OL��F��.`A�K�t ACROx��Q1��ND_C���i��A�d��ROUP���R_�н�E �Q1 �h�s��y���y����x
��y��y$�hAx��n���AVED�w�X��ueQs:h $���P_D�H Y�^RrPRM_��1_HTTP_i�Hx�wi (*�OBJ��l�b��$2�LE�3��P���j � (#��L�_
�Tp#��qS�P�c��KRL{i?HITCOU��3!6�L`��Q��U�`��`SS��J�QUERY_FLA�r�HWR�N1x��kpgPINCP	U����O����Œ�!tƑ/tƑ��IwOLNw�l 8!�yRu�X�$SLL�$INPUT_&Y$;`�P,��M �SLY�x�m���M�I��C��B��{IO��F_AShn}�$L��Ӈ��8A�b_1���V���@HY1�̡��NqUOPeo ` ���2��¼���æ�[`P�c;`
�.�æ;��$�s�UJa�p � K�NEaG4�v72k�Da��2J7�s��+J8��7�I_1��>��7_LAB�1�Px��ɸ��APHI���Q���D�J7�J8*é_KEY�� �KǐLwMONx�q <���XR����X�WAT�CH_��C��i�E�LD��y���er� @Р1V�wFP{�C�TRCz��%�L}G��s� !�/$LG�Z�R�`��c�ƈ���FD��I����\!���ȍ �� ��e�Dqf�ce���e� ��e�� e���@0J�_�ѐ1�ѫ�ژF �A�׷���Cd(��SB����c�ֈ�������I���؅��֘� ����RS=��0 7 (�LN��<t��7���N�	�D[��U��i��PLr�nh�DAU��EA��0h��T���GH�R4�BOO ru�3 C���`IT������ ��REC��SCR��#���DQ��r�qMARGX~p#�,����dM�>�����Wp+���}䟣JGM���MNCH�s��FNt�K��PRG���UF��b@��FWDv��HL��STP���V��� �����RS"'	HzP����CdD 1R���_��	U����@^���m�������G��@PO�

���f��OC/ ��EX���TUI��I#�\� 7h�Bt�B���<@@<���e��<@�N�q��3ANA��A2x@V�AIɰ�tCLEA�R�FDCS_HIP$�!s�O�O��SI��S�B�I�GN��<��é�T܅t�DEVaLL�Q��_BUFF�	1vu�j@T��$��EM������V�*A�bwu�j@����zq�POS1�%2��%3�!c���
0x �h��x�Q@5���.�IDX�TP~B?baO� ��1"6ST��R��YmrD1 w$ES6CS;����b6u6���#��_�y L����`Ϩ����`Na�eE�p�e��e��?_ z ��\�𢀣r�C�MC�\�{ �h�CL�DP�UTRQL�I��Ty�8I&DFLAGmr&@�QZC�Di��ZG��LDZEDDZEORGy�]mB�ظq�` ��D!s�D/r C|�| �G�DD^5DZE�S�PT8@`��@T>VRCLMC)T�O��O;Y3��A���_�}�'�$DEBUG|Gu��XDATA~�r=�T�@�UFE��=TmqC�MI6p^�g~ de��!RQo�=G�DSTB�`0c �V;��XAX-B���WlEXCESH���"�RMZ`^�S 	�R-D�}��RSq_�����V_�P�X��xk
oh_�MJPTmā K`������aMICb� � ��0�"]w�R+CT �NS��fR���gA�jL�bC�`C�s��aUSED� O�� ��CURPXk_T�Ql�PS�� �A|�NpTtZER�p�pyS�`E�B_FR(P��8q�vZ_�Ѓt���l�A�PAKmă �\����6�UB��L�IÁ�sREQUI[RElMO�|O�{��RB�@L�0Mlń ��������s)R��MNDz�S�"�c�Z��^�D���v�IN���v�RCSM��x� �a�1�E�D��AL�PST�+� � 4)�L�O�`�$RI% �%EX��ANG�"�Q8a�ODAQlŇ�P1$ql��MF��� &�9�2� �5K�W��V�SUP�5YaFEpR�IGG�� � �fP�3VѲS�3v�4I�ΰ%C3������������`���Q'�PET!I^�� �aW�M��^"�� t�MD�I���)��)�iQ&�H8􀚱)�DIAͱ*�ANSWQ�)��!:)�D��),�\�\P_�� �aU���Vg�\@�QAOD�_{P^� �h�3�L}P�}��ڨPڮh2 ���P٨KExF���-$B��ͦ�0�ND2kRB�*�2_{TX�4XTRA�4V����LO��_�1�Ibl��R�k��R፡�������RR2>�U�0 #|����AQ d$CA�LI�PW�G�ȷ2�� RIN��̳<$RְSW0GT��wABC$�D_J<���qϰ�_J31�
�+�1SP����ϰP�+�R�3Qͦ�d�ϰB��J����BQO]!�IM�dRCSKP GJ�ģ�~���J��dR�Q�����������_cAZR��#�ELB!<��kQOCMP��eQ�71n�RT�QN�~�11���l�01�p�c:~�Z|�SMGA �vbTJG�0SCL,`�SPH_�dP�����B�ϰӰRTE�R�̳ �IN��AC�"�����E�X�Q�Ң0_N��� �@�$1dQ� �db�%�cDI9�eP��DH,`tX����� $Vհw���c$��怳A(� �"B��`R������H �$BE�L4�d���_ACCEL�������`S_R��Q �aT71Z#3OqEX+BL[r �@C����s��Sq��h>���>�3[sRO/a_�!��o�u�R�*p���_MG!$D�D�����$FW��P���������D}E��PPABN�RO��EE��!���8@���!~Q�P��[pR1q_԰~P�`C� �~Y���Q �1YN�PA��\��@�\aM�Q�����OL�t�INC��������R����QENCS�԰��R����TPpI�N+2I[r����N�TVE� ̳23�_U���" LOWL�H k�8@�@DF�T�P���0��b9C�MOS  �d��`u�WcSPERC�H  ]Otp��  ����ʑCbTʑIאA�FNr��A[r�L <�Ùg��k�C>&�YTRK��(1AY ��Mstan![r}%r#�pT�xa�80MOM����Rtb�@���T��ȷ0�#@�!��DU��\r�S_BCKLSH_C[r 5�P~tpd���4�):s��CLALM�A� d`[5�CHK8@�04�GLRTYΐ�����Ar�_@�s_UM�S��6C�S����3 LMTN�_L�@<��4P��7E�=@�;�0�� E��c��S"FD�P	C��Hn� ����5�C7P]����CN_b�NGS�F�SF���VF�1���zA[r��E~HCAT�>SH @�㲤��dq�!�}�0\q}�qГ�PA�4�_P�5�#_����u& ����#�T�5JfqB`̋S.OG�G�"TORQU8 f�q�)��`�r��!���R_W�% n$zѓ�d��e��eUI"kI0kI��F�``a��oh����VC��0)�$�c1�n��o���fJRK�l�b�f�, DB��Mң, M�u�_DL��"GR�V!dt��t���aH�_���cA�HzCOSU{V�UxLN�`x{�e t��zy��zyLa�z�|�ja�eZsp��aMY��q�xar#�i{�TH�ET0INK23���?�~�pCBD�C5B~�CذAS��i�`Ldw���w�D�SB�㜕�O�GTS��C�U��t�`S��ˊ�s$DU�0"'��Ȳ��b ����!QʒZC�!NE��\�I�p�3`�0�$b�3�A7�`�i�8GuRxRqLPHUu>�>�S�e���u���u@>��vۓŚ�vb�V��QVw�t���V��V��UVěVқV��V�V��H��$�����QT����HěHқH��UH�H��Os�O���O-���O��O��O�ěOқO��O�O�vF>�d����uŴu��SPBALANC�E��bALE��H_7�SP�ѕv¤v�>�vPFULC�C°+�C³u�1�P�U�TO_�0�UT1T2����2Ng1�� �īѨ!E�#����!�T/ O9���`IN�SEG��bREV8��bDIFX%*�1��V�1�K O!B�K1$s�'2�P�r1tLCHWAR���y�ABgQ�%$MECHm��{���6AX{!P)D��Y�e�y�� 
���Q��n�ROB�CR�R��ՏB|0�MSK_|���� P ��_6 R����Z$1�B�)4��c�IN���MT�COM_C�`����  ������$NOREv���S�e�� 4� G�R�R��FLA��$XYZ_DAv��3 "�DEBU���X��S��� �$TwCOD:1 ����"��� $BUFINDX <����MOR�� H �� ��j6!� �)4Ҹ��A5��0{TA IB_����"G� � ?$SIMUL�P��������OBJE|���ADJUS�����AY_I�Q�D��OUT�P��� � �_FI�=�T 
`������7Ж ������ ��DQ FRiI37T5RO�P�� Ea: �OPW�O�`��,��S�YSBUP��SO!Py��`1�
U���PRUNU�PAB"�D�����_��-B� 7�AB��/@��/IMAG:1�&��P��IM8�IN�p� RGOVR!D,����P� ����L_w��QM�2��@RB@# ?AMOC_ED��� /@�NP�M|.A� MY�19-A���,S�L��� ���OwVSL��SDIZ DEX�C��C/!�	V`�N��Q� ������#C�@T�'!��_SE9T�P�� @� F"�� 1RI����\#_q�e'~!q!Z�ѝ�.�@ ��T�ЪP�ATUS� $T�RC(�' �#BTIM�'�!I��4-A��#z�� D�E� ��"Y�Eҷ!��8  K0�!EXE� �1 q2%2�$N#�U �Ƽ UP��415 ISXNN�'�A��a^�)L�PGc�q $SUB�!��{!��!#JMPWAI2PP��5LO	@�������$RCVFAIL_C'� �1R ���ӊA�@�D�мE�pR_PL#D�BTB�Q�B� BW�DF~�UM�P
DI�G���PTNLP
DeBRLy�P�P<�pPEEDZ0�CHADOW�P��~��E��D��1DE�FSP�� � L���@_�@���C�UNI��'�@h1R�,02#L ���P�!&�P�PV�����P@��� ����N4�GKET&R`��.P�PYB� h ߀SIZE�P�� ���QS��OR#F�ORMATp�ODC�O��Q��EM����T	SUXh �B!PsLIJB� $n�OMP_SWIT�J�E��W��o�Z��AX/@J@AL_ C��P�@G��`Bo�i�C:�D�$E�41�J3Dh�{ T{PPDCKh|���CO_J3���8bvb�;�.o@m��"`C_TAf �; ���PAY�:��d_1�j2�c`J�3���k�ev�c[TWIA4y5y6:�MOM2�)sIs6sIs4Cs`�B�0AD)smv�6smvCsPUx�NR Nt�u6s�uCr�2�Q���` I$PI 5��e��eO��e���e ���ez��������������1�ђ�_%�CHIGc�C�5 �D���D�5@ ��ă���A��A�5SAM��$� �����5MO	V��I�L�/��N� J�>��H��@�`W��`�J�U Z&pF�`H��H�IN��`䃖� �����2��ؘ��؛���GAMM춿!���$GET�D��dT�
��LIBRt^1|BI��$HI]0!_� J�m�EG�z�1At�����LWo��� ����٦���b��r@!a�C@EU�:�  dnI_�W T�b �ha~�B�IsT�mvA��c �$Qh W1���I} R���D;�c�f1�4e�LE@E��!θ�h���@_MSWFLDM`SCRn87���N���y2�@�QA��P��UR	�I���p�S_SAVE_DXRg�`3NO�`C�! a2�dg�K��o�q�i| 
��i"�����@��bH���cD���H��@>� e�Q�I㈈~���Ĉ@e�a��A�a1hRL���� � G�YQL�s��~�=�S�� [U��%@����o��� ��	�.��W���A�p�V��M�#�CL"�q���%��1y2�PMX�O"� ό $��l$Ww�6���aw��d u�du�du�Cd0@4��P��S``XPO��caZ���P��z�[ ���OMp��f��ϻ�������:pCOIN��4��R�a_�2� |ba1�g�Iy�� 6s��Csg�"z����<z@aE�)P�r��>®)P��`��P�Q�PM��QU� � =8:PQCOUr�� 7QTHT@HO��l 7HYS�PES5�k�UEW ]�jPO�T��  �PPU�e��"U�N� ���{�� P��5I�3|B�ROGRA�!��224O �ITİޙ INFO}� ��Q�
)���r�O�I,� (M�SLEQ�Ts�T�-P�OS��4� 4�:PENAB�� PTION#�DM��\�D�GCF��U"�J@a��Q�R������OS_sED�0� �s R��KA�_#l�E��sNU>'8(AUT��;%COPYA�]0\,�A��Ms�Nf j+��PRUT�� m"N��OU b�0RG�ADJ}�yRX_���B$P�&��&W�(P�(ܰ�&�C� ��3EX @YC��^�RGNS������LGO �@`NY�Q_FREQ�rW`�r�r1�T�LAĳ�i1�!Ds�eCRE�X�w!�IF��NmA	�%�4_G�D�TATg@�4c�MAIL�W��1аg!Qx�1V�D4ELEM�� ��@�FEASI�e�4�q���)B@ep�[F"{�W�I�U�i2j�o2 ӳ�BAIBaA`E� ��VA�FBASKb�EW��qqU��� |�$�A~�GRMS_TR�C a���C�㸀��A�D� C5����	~gB 2� �� �䬔MV�BLWRT�������BxW�wȴDOUd���N�F2PR��z��[GRIDއBARS�TYȟ�z�Odp}� �_�4!0�R�T�O���� � �POR�c�v.bSRV�0)<d4fDI��T�`Uahd1��rgh�rg4pi5pi6Jpi7pi8Ta��F(����� $VAL!U�CZ�MD)�a��� �~��bc�1W� ANY���b�1R( w1W�TO�TAL��qWsPW�_3I�QmtREGENkz�rX�H�w53"vR TR�C��kqC_S]��w�p#V�!
$�r��BEC�PqpVҵR 4sV_H�P�DAR��p2�S_Yh����6S,�ARR��2� �"IG_CSEh�p4bE_� F�C_�V�a�U��p�_lF�{��SLGj�
���c5��T�dUp^pS��DDESaaUc����ހTE��>	p�� !�q0���qJ����=CIL_�M�4`�ѳ�p�TQ@R [��@���V��EC��P9�HA��M��[V1��V1ɛ2؛U2ɛ3؛3ɛ4؛4ɚI��p��J�1�U����9�INf�VIB�b�����Dщ�2��2���3��3��4��4���}�|Rہg����D $MC_F,u "�J�Lh�g��"HsM��I���S� ��[��q�K�EEP_HNADED�!H��@R�C$��0h��Q���i�O KG�� �X�i��1�3.i�REM��h�]qPb������U�4eh��HPWD  �H�SBMSKbCOLLABT�pe�4Iq�2DITI0�ซ!��� ,M�F1L��|�r�YN��V��M�C���lpUP�_DLY}�ŤDGELA��^q�2Y2 �ADR��aQSK;IP��� �,`� �O��NT^��Ѳ�P_� ���� ����� �q�Ɋ!�ɉ`�ʖ`�� �`�ʰ`�ʽ`���`��=9	1�J2R)0�ǖX�@Tl3�� '���#@D���D���wRDCx�� ���ER�RV ��n�R�1p��o��OTRGE�8yC�ӫRFLGL��$OTSPC11U�M_��F�2TH2�N�Qa��� 1�� ��P! 11�� l��$�t��,�AT���#S��  v6��� ���! OT�ℽn�H�����z�2��ʈ��������@0z�3�����)��;�M�_� z�4��̂�����������
��5�����#5\GY z�6���|����� +z�7����0/AS ��|�8���v��������S�q�  Q{�p,��㾰-EJ4ҥ�;��"LNv�#IOC��)I1 ��ar�POWEh�G� r U������Ht �P��"$D�SB�0�0BGs��C(g��"��M/U�P�)�D� PE�2ǐM�DG7��M!e� D���7DBG_�PP0�TSJ1�qPG/QAP���3��S232N�%� ����u��ICEU�BFp�4���ARIT4�FqO�PB4�&�FLOWc�TRM Srͱ�P'��CU�0MJCUXT�A�'�INTER�FAC�4��UBp�eSCH3Q� �t9��G1��6�$L��OML��A�"PI��@vPAP�� 	Ti Cc�p���H�C=�EFA"�@�=�:���c� ���p]r Ė��b m��F0Q ���"Ł  2� ��S��r�	�' �$N���U�/u�7SWp_J�BVDSP�NVJOG�p�3��_P��BON�К����L�.FK�@_MIR�jQ�4��MT~��SA�Pp���Y��P�DGQS�?��P&�GQ�0�UBR�KHaA�Fb��b�� bʃb9RP�@$�7S��PBSOCBV��N�>eDV�Y16"��$SV��DE_O�Pl�FSPD_OKVR4����Dyb&|SOR�g Np�f�F`�ggPOVjUS!F�j���cQ�F�fE��L�UFRA�jTO�DLCH��W�OVxd �gPWv��gS��E�K`vP��  �@;�TIN��1/$OFShpC�@e�WD�a+t�aJa"�U�d`TRA�2�QFyDг�QMB_C:�
�rBZPBa��F��r�q�SV��q��@��d�ùbG�w�XAMC��B_b@�Rr-�_M��p'B3��"_pT$C�A]P3�Dbd�HcBK�A�Fy�IO %q���!��PPA|����������8��"_rDVC_|0w3ꀤA2 ���a�͠�R��3	�Xp�u�7@�PxaqUw3\P�&CAB�Ѐ"Q��pÿp�^�O� �UX�FSUBCPU 2tPS��� г �t�@Ѻ��s�t�"��?$HW_C���@ї��� ��'�$U3�d��ATTRI�@"�tP�CYCL��NEC�AN��SFLTR_2_FI2#9T�6v8�LP�[CHK��o_SCT�SF_�cF_���*�FS1�r�CHA�щ��8�rB�RSDz�10+a�C1� _T�~��:��s@EMG ��M"cTϢ��Ϣ���W�DIAG�ERAOILAC����M��CLO.`\�Tf2�"�bX� ��X�$�PR�MSP� ^@��C݁z�0	QsFUNC�6ARIN�;�$0i��A��S_GPO d�	���r�	�#�r�GCBL���:�A3�/�6�/�DA`
�t�:�3�LD�@l`����dOQ�����TI�����2Q�$CE_gRIA4�2AF��aP�3��Jp��T2��1C�C
��qOI��vDF_L~ r�A�@�LM�3FAE0HRgDYO�QrpRG���H��a |�;�MULSE+ЦC��]`�$J�jJ�b�g�k�FAN_ALML�VC��WRN��H�ARD`�F0��2$SHADOW%p �0��v���1q�UY_&p��AU֠RԤ~(BTO_SBR�$�D�[PM��߃�e�M/PINF]p$�x䜒���REG!&��D�G��p�V�@#fDoAL_N�tFL �^�$M������0�tpq�p $2!3$YM2{A R*3��� ��SE!G� 7Sl`/�A'0�$�Te2]c>�`��UAX�EQWROBNZREMDNVWRE0a_���0cSY	`i�`��S���WRIE0B��SAT� OS)@`�`E�AD K���%�GPB���^q5��>�OTOr��D JpARYNS`8��>���PFI�P~�S$LINK*��GTHW�@T_���^qJ�6^b�X�YZ�B�
7�OF�FfpW50� s� O	BLPղ�;q@�@�FI=��7@3ddղfT_J�1�B�b d���8^b�0� �.y�fC� �VD�U|rI�9��TURB��X�ßFs�X���0NFL� pm�<����30^btq W1�D KsPM��Te3Ƒ��������|CORQ2�[Q��֑���PO��N��m%�C8YQ��$OVE�!M2MU@o!�%	�%�&kA�'o��'��$AN�Z�!��N1�!�P � &��!�%�!�',5	�,5�#[QERxQ�	B��E-0�p��j4A1���-�D{�x�{�AX;s�B{�>��� Y�5]��9���9���: ( �:� �:� �:_�:��:1��6;��9;� �9;��9;��9;�I;� I;�,I;�<I;�LIiA�]IDEBU�$����U�Q{r{AB�{�y��a�#Vn�� 
(R��PU֑\W ]a\W��\W(\W�\W �\W_\W���k��\Y�LAB�N%��GROg�N��W�B_;�Q6���c � J�f9aO%5e8�AfAND ��_4X��b18�~g W����h0=��hZ�� NT��/s�`VELA��$�ay�~�f�SERVE�`N�� $� �Aq!pPOmr�p�2 	q��b1���  $&rTREQp�
%s��/p�3w���2�Du��v�_ �� l˰�q�ERR�2I��`�$N�qTOQ�$� Lm�P�4��v-�Gu%m⋢�$t��.q� ,h qHubp�1RA�q? 2� d	���q��r;p ����$� @�о2�d_�OCl�-��  }�{COUNT���!��FZN_CFG.q� 4됺�`�T��'�Sɐ���r�$py��� �MPM㠔��H��#�!���FA��	5���X������q�x�t�t���Po�$pHE�L��~�� }5��B_BAS���RSR��ɰ��SH���r�1�wr�2��U3��4��5��6���7��8�we�ROO0=��p^ � NL	�q�ABss�s�ACK�9VIN7�T����$�U�r�ԡ%�_PUX{��Ї�OU=�P����R��vՠ��6TPFWD_KAR�qL��pREtQ�PT ���QUE��-�� z����I��<SR��� ���`��SEM�XQ�fQm�A܁ST�Y4�SO�.�DI�@��ࡩ7�_T}M��MANRQq�� END$$K�EYSWITCH�����S��HEzBoEATM �PE?�CLE�r�!`ɸU���F���SX�DO_�HOM��O��(�EFf0PR��������A�C�O]шp�qO�V_M@���IO#CMl�d!CrS�;HK�� D}����U�ޢM7𲤵 �mFORC��WA�RM�!�S�OM@� �� @T=�U���PX�1��2��3���4b�E�<�O��L�����r��UNLO�^��3�ED� � �SNPX_;AS�� 0���|�� �$SIZ���$VA?`�uMU/LTIP�S����A��� � A$m�T��� g�S���'�C�p��FRIF��27�SȠ��ķ�N=Ft�ODBU��``����u\`�Ss�n�� xzpSI�r�TE�]"�SGLO�Tf�&��h�c<��P�STMT���P+���BW� Q�S�HOW��0�SV�\0_GĂ� _$�PC`8�\3�1FBZ��P��SP�A?����EpVD��Â��� �|qA00 �d���#���#��#�T�#�5!�6!�7!�U8!�9!�A!�B!�@��#��Q$�#�F!��\@��-�1:�1G�1�T�1a�1n�1{�1���1��1��1��1���1��1��1��2� �2-�2:�2G�2*T�2a�2n�2{�^T���2��2��2��2��2��2����P-�c �G�3T�3a�U3n�3{�3��3��U3��3��3��3��U3��3��4�4-�U4:�4G�4T�4a�U4n�4{�4��4��U4��4��4��4��U4��4��5�5-�U5:�5G�5T�5a�U5n�5{�5��5��U5��5��5��5��U5��5��6�6-�U6:�6G�6T�6a�U6n�6{�6��6��U6��6��6��6��U6��6��7�7-�U7:�7G�7T�7a�U7n�7{�7��7��U7��7��7��7��e7��7����VPǰ=U,r� 5p�P���
����a�z��8`RѡCM���rMbpR^pE��dQ_P��R�`�uMq���cY��SYSL�p�`� � q�'⏇��f����`0��"d��VALAU��J����Q[hFa�ID_L�eHI�~jI��$FILE1_q��d��$�:��cSA+�� h�  �VE_BL�CKˣ�bj��hD_CPU yr� yfК�ȱo�d�pYO�k�R �� � PW�R���aqLA���S*�fswqptRUN_FLG�uet�qpt@���u�qet�qpuHk��|t�ppt�TBC2���� � (�B �pM���;�� ��.�'TDC�p��!�π��/��TH.�J��T�V�R�4�ESERCVE!�w�.�w�3t���$$CLAk� o���P��OЍO� ���զ�����׹�I�RTUAL����A�AVM_WRK �2 �� 0  �5����'��J� J��]���O��!�o�������]�Н�ܟl���)�1���B�S��� 1Ɖ�? <�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f��x��A�C1�AXL�MTÀ���Z�  d��IN����PRE_EXE��1����QAT��R�����IOCNV_�NUM�� ȶ�P��US��V�@�IO�_$� 1�P $�痑�����?����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v������LARMRECOV ������[�LMDG �k�v��LM_IF k����5� G�Y�k�y�#��������ҿ�, 
  �χ���2�D�V�h����ANGTOL � � 	 A�   �Ϲ˟�PP�LICATIONg ?�������ArcTo�ol �� 
V�9.00P/03���y�
8834�0���F07�$�1�612������7DC3�y���N�oney�FR=Ay� 6Tݚ�P_ACTIVJ������UTO�MOD
����P�_CHGAPON�L� �OUP�LED 1k��� Y�]�o����CUREQ 1k�W  T�������	�������Ф���_ARC �Wel��AW����AWTOPK7�HKY����� ���Q�c�u������� ��������)� M_q����� ��%I[ m������� �/!/{/E/W/i/�/ �/�/�/�/�/�/�/? ?w?A?S?e?�?�?�? �?�?�?�?�?OOsO =OOOaOO�O�O�O�O �O�O�O__o_9_K_ ]_{_�_�_�_�_�_�_ �_�_oko5oGoYowo }o�o�o�o�o�o�o�o g1CUsy� ������	�c� -�?�Q�o�u�������0��Ϗ	��TO�������DO_CLEA�N)���`�NM  ��������П������_DSPDR3YRg�:�HI���@��b�t��������� ί����(�:���MAX��G� ��8�X�XG��T����PLUGGG�H�T�X�WPRC�B����Q�C���O��"���SEGF �B� �� �����b�tφϘϪ���LAP?�R�� ����(�:�L�^�p���ߔߦ߸��߿�TO�TALz���USE+NU?�L� -�1����RGDISPWMMCB�J�C�O�@@��L�O=��_�-�RG_STRING 1�
�M�S���
��_ITE;M1��  n���� ����	��-�?�Q�c� u����������������)I/O SIGNAL���Tryout� mode��I�npi Simul�ated��Ou�t{OVER�R<� = 100���In cyc�lo��Prog� Abor���~estatus��� cess Fa�ult�Aler��	Heartb�ea�KHand? Broke>; =Oas�����C���C���� ///A/S/e/w/�/�/ �/�/�/�/�/??+?p=?O?a?�WOR� ��1/s?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O_^PO��=P�;&_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono��o�o�o�o8RDEV @^�`T_�o,> Pbt����� ����(�:�L�^�PALT����? _�����я����� +�=�O�a�s�������ໟ͟ߟ�s�GRI ]���)����Q�c�u� ��������ϯ��� �)�;�M�_�q�������R�ͱA����� ��+�=�O�a�sυ� �ϩϻ���������x'�9߻�PREG�� r��Kߙ߽߫����� ����)�;�M�_�q��������?��$ARG_�0D �?	��� ���  w	$?	[4��]4��?U��SB�N_CONFIG� �srm�C�II_SAVE � ?����T�CELLSETU�P 
 �%  ?OME_IO??%MOV_H������REPм:�UTOBACK��� ���FRA;:\_� A_֖��'`� _׊� ��� �23/04/0�8 11:47:14_�V�_��	6-{��V}� ����_քk/ /)/;/M/_/��/�/ �/�/�/�/�/z/?%? 7?I?[?m?�/�?�?�?��?�?�?�?۰�  �v_Y_\ATB�CKCTL.TM�P DATE.D���DOVOhOzO�OSIKNI�����S?MESSAG��A���(�KODE_D ��������EO�`�O�SPAUS=Q!�� � ,,		��  �M_[WA_ {_e_�_�_�_�_�_�_ �_�_/ooSo=oOo�o��� T*PTSK � 0]��OV UP3DT�@�Gd�`�F�XWZD_ENB8�D��vSTA�E ���e�WEPLSC�H Rb   �fj|�� �������0� B�T�f�x��������� ҏ�����,�>�P�nDsROD,r2 ���Lڳ�� %��ɟ۟����#� 5�G�Y�k�}�������WEROBGRPƮh[r�b��WEWELn�������� ?�Q�c�u����������Ͽ����
�XI-Ss�UN� ����ա� 	 ��E� ��������eI�_�T����pϩ�T�Ϧ�:����	���ϻ���.��1�METER 2�f�� P�t�����+�SCRDCFoG 1 �l' ��������߀��'�9�K���Q ���ߛ��������� \����=�O�a�s���`����8�KYGR;���`_��@NAME7 	�	Y���_ED�@1��� 
 �%-%@EDT-��#�Tx��� *�? G|ځ0��'�?������2�"�6�G� �}��l��3�%/I[�I/ ��8/��4�/� �//[�/?\/n/?�/�5M?�/�?�/[�v?�?(?:?�?^?�6 O�?fO�?[BO�O�?O�O*O�7�OUO2_ yO[_y_�O�Oh_�OB�8�_Y�_}�\��_Eo�_�_4o�_�9}o�_�oo�\�o`Xojo �o�CR�  _��V]p�"4��X��# NO_D�EL����GE_U�NUSE����IG�ALLOW 1��   (�*SYSTEM*��	$SERV_�á|ٕ�POSRE�G��$��|ܕ�N�UMÊ�֍PMyUA��LAYM��|�PMPA�LT�CYC10�"�5��#�[�UL�SU�׍7�����Lq���BOXOR=IǅCUR_��֍�PMCNV����10K���T4�DLIB����	*�PROGRA��?PG_MI#�M�F_�AL-�l�V�_��B����$FLU?I_RESU;�ï͏�s�|��"� 4�F�X�j�|������� Ŀֿ�����0�B� T�f�xϊϜϮ����� ������,�>�P߳x���LAL_OUT� �����WD_ABOR<�e����ITR_RTN � �d�����NO�NSTO �� �M�CCG_CON?FIG 
�����:ㆃD�R��E_�RIA_Ib����z����FCF�G 
.��mރ�_LIM��2�- <�� 	������b<���-����`���PA��GPw 1���A��i�{���L�C�������C1��9��@����C��CV��]*��d��l��s��d��C[��m��v���������� �C���D ��g?��HE����]�G_Pݐ15� -�P������\�HKPA�US��1��z� K�(n��\�� ����/�*// :/`/F/�/�/|/�/X�O�����g��COLLECT_��a��М�7EN-�p����2�!NDE3���P��r1�234567890o7�b����m?6�c'
 Hy��c)�?�? �|�?�?$O�{�?OhO 3OEOWO�O{O�O�O�O �O�O�O@___/_�_ S_e_w_�_�_�_�_o��_�_o`o+oI6���; ��I6IO !X91�h���o��o�gTR0�2%"�m(�`�i
Ao&~�"�#�mPzn�i_�MOR��$5� � R	�u���y�����9�'��r+��%�},�n?WW����`KT���aZR��&�/�ŏāĂC4  A�����`x�`A���Cz  B�C�0BO 	�C  �@���`�a:Wd�
��IQ3'��}��T_DEFx� l�%^y��M�INUS:�mz厔�KEY_TBL � 4�z�Ā �	�
�� !�"#$%&'()�*+,-./x7:�;<=>?@AB�CP�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������S����͓���������������������������������耇���������������������a��LCK��鲐���STA�ߌ�_AU_TO_DO�����IND04 �1Rg_T1��T2Z��� �A���XC*� �2(���08
S�ONY XC-5�6ɏÁࣀ�@����1� Kp�w�̵HR5�98Ns���R57�"�Aff.�h��ϖ� rϻ��Ϩ������ '�9��]�o�Jߓߥ�p������i|TRLO��LETEo�J�T�_SCREEN �5�kcs�c\U��MMEN�U 1)5�  <��g���^� ���#���������� /���e�<�N�t��� ������������ (a8J�n�� �����K" 4�Xj���� ���5///D/}/ T/f/�/�/�/�/�/�/ �/1???g?>?P?�? t?�?�?�?�?�?O�? OQO(O:O`O�OpO�O �O�O�O_�O�O_M_�$_6_�_ylA�_MA�NUAL��Q�DB�wq~r��DBG_oERRLU�*M��a �_o*o<n��QNUMLIM���`d��,�DB�PXWORK 1+M�o�o�o�o�o|�og}DBTB_��G ,�]؃HqÄ��QDB_AWA�Y�S�GCP μ�=��lb:r_A!LX` �6r�RY��	�t���X_�P 1-��+q|�
�o��Ȅ���h_M7�I�S��E{@���ON�TIM����ɼ,��y
���sMO�TNEND���tR�ECORD 13�M� ���sG�O����{Er� � �$���,�S�w�� ������V�l���d�� ��=�O�a�s����� ��*�߯�����9� ��]�̯��������&� ۿJ���n�#�5�G�Y� ȿ}�쿈�������� ��j�ߎ�߲�g�y� �ߝ���߬ߺ���f�f�-�?��c�N��� ���p�U������[� ��4����wt�g�y����������B��|DJ_��-��Q< J�����>��TOLERENC�CtBȌrQpL����PCSS_CNS�TCY 24zi��P��r�DRd v������� //*/</N/d/r/�/��/DEVICEw 25/ v �/�/??1?C?U?g?�y?�?�?� HND�GD 6/#pC}z�>LS 27�-�?O-O?OQOcOuO��O�?!PARAM� 8�ysr�U�D�SLAVE �9�=�7_CFG �:�O�CdM�C:\!L%04�d.CSV�O�pc�8_�RyA eSCHmP�1��Nx_�_�G��F�R�Q�_�Y�QPJP��S�^�q�q�LRC_OU�T ;�-q�O_?SGN <�������mE15�-APR-23 �11:34hPQ708�h48hP�& V�^�i�a�N�`ya@�S�Þ�j��a��n�CVERSIO�N ljV�4.0.1 �EF�LOGIC 1=^/ 	�XP�Py�Q`}2rPROG�_ENBw��6�sU�LS7� �62r_�ACCLIM8����C��sWRSTJN��偃Q�2qMO�|�Q�B �I?NIT >/��vQ �vOPT�@� ?	=��
 ?	R575�Cj��74o�6p�7p�50��%t��2p��X��|,wM�TO  Y���o�-vV$�DEX��wdtb`+�PA�TH AljA�\�x����HCP�_CLNTID y?v�C k��ʟ�IAG_G�RP 2C
Y ��� 	 �D�  D�� �D  B��ff���?����<��h�V����B�N�C�-Bz��Bp�e`��mp�2m7 7890?123456������  Ao��mAj1Ad�A]�
AW�|�AP�AJ�-AC/A;��A4-�ؠa@ɠeT��A�A�hPB4���� ��Y�a
עu���ApffAj��yAeK�A_�AY��ASy��MC�AF��A@ �9��"�4�9�xH�9�W�@�X��ȑ�@��y�������ſ׿鸃;�d5?@~f�f@x1'@q���@kC�@d��D@]��@Vv���-�?�Q�c��s���l��@e�@^��@W\)�@O��@pP@?�!�7K�@.V��Ϲ��������S�@M�G!�A���@<1@5���@/l�@(�w�@!���\3� E�W�i�{�]��/�A� �e�w��K���� ��������=�O�-� s������A���x������Ѩ�/�>���R��?�33?Y�������/�7�'Ŭ6 4��F#��L/�@��p�?�
=@�@�Q�OZ�m@,�AheP�eP��9�= c<���]>*�H>�V>�3�>����/�<���<�� ���^ ��?� �C�  �<(�U�R 4;�33����	��A@�R?7���)�� 7]o;��{�?�����/��?��73!>�(�>���?!=���/��7�G�[/G�/��Ґ�Ռ%����eP� @����@hP@Q��?L��������Iߟ5�˦�G?�"��'�p%10?{&���L4V?5�C�qP�̇�C'^?�,�?�? 7<�P �?�?��?�T�?O�?=O�+r[HgH�DD@Ob�Dq�C3���*�?³��@F�/O�O+O�O�O�O�O_�DIC�T_CONFIG� D����d�eg�U�ST�BF_TTS�w
@�ywSp�s�Q�V/`�MAU�p��rMS�W_CFKPE�� � �lOCVIE�W�PF�]:��� ޟ0oBoTofoxo�o� o�o�o�o�o�o�o 1CUgy�� ����	���?� Q�c�u�����(���Ϗ ������;�M�_� q�������6�˟ݟ� ��%���I�[�m��X�����\RC�SGg��R!?���ۯ���4��#�X�G�|��TSBL�_FAULT �HΪ�X��GPMS�K�W��?PTDIAOG IOY�A�)�UD1: 6�789012345�\X=P_B�T� f�xϊϜϮ������� ����,�>�P�b��8# t:
1Ϫ�>9VTRECP߿�
����?*�'�9�K� ]�o��������� �����#�5�G��߀���ߏ�2]UMP_OPTION�P����TR�R�S����P�MEU��Y_TE�MP  È�g3BȤP$ �A! UNI�P�U$Ѷ�YN_BRK �J	o<REDIT_~��ENT 1KΩ�  ,&M�AIN_MANIPULAC��P���P&DESCA�RGA_INDE�X� O�\S&C�APTURAEQV�EY� ��CL�_�CO�'�L�_��%�	IR�_A_HOME yXW��&P� �E���
PIC;K_w RAD�.�
����l�,/\R�/W/>/{/b/�/ �/�/�/�/�/?�//? ?S?e?L?�?p?�?�?�?�?�5m MGDI_STA7�Q$�R�m NCC1L�[ C�[�MO@O��
��d���O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o ��8oJo\ono|i�A|o �o�o�o�o�o�o  2DVhz��� ����
��j1o;� M�_�q��o������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���)�3�E�W�i��� ������ïկ���� �/�A�S�e�w����� ����ѿ����!�� =�O�a�{�qϗϩϻ� ��������'�9�K� ]�o߁ߓߥ߷����� �����+�5�G�Y�� �Ϗ����������� ��1�C�U�g�y��� �������������#� -?Qc}��� ����); M_q����� ��/%/7/I/[/ u/�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?/ O/OAOSOm/_O�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_O�_'o9oKo eOwO�o�o�o�o�o�o �o�o#5GYk }������o o�1�C�U�ooy��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ�[���)�;� M�g�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ��!�3�E�_�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿����������+� =�W�M�s����� ��������'�9�K� ]�o������������� ���#5��a�k }������� 1CUgy� ��������	// -/?/Yc/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�OO%O7OQ/[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�?�_o o/oIO;oeowo�o�o �o�o�o�o�o+ =Oas���� ��_���'�AoSo ]�o���������ɏۏ ����#�5�G�Y�k� }�������ş���� ��1�K�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��7�����)�C� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������ ���!�;�E�W�i�{� ������������� �/�A�S�e�w����� ����������3� )Oas���� ���'9K ]o�������� ��/�=G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?���?�?	OO 5/?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�? �_�_oo-O7oIo[o moo�o�o�o�o�o�o �o!3EWi{ ����_���� %o�A�S�e�w����� ����я�����+� =�O�a�s�������� ��ߟ���/�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������͟׿��� �'�1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ�� ſ��������)�;� M�_�q������� ������%�7�I�[� m�������������� ���!3EWi{ ������� /ASew�� ������/+/ =/O/a/s/�/�/�/�/ �/�/�/??'?9?K?�]?o?�?�?� �$�ENETMODE� 1M%_�  �����?�;�0RRO�R_PROG �%�:%�/O<I
ETABLE  �;�/{O�O�O�G
BSEV_NUM �2  ��1��@
A_AUTO_?ENB  �5�3�D_NO�A N��;�1�B  *U�'P�'P�'P�'P��@+&P@_R_d_ TH�IS�C��0�K_A�LM 1O�; e��'\�+e_��_�_oo)o;oi__\�BP  �;%Q��2�j�0TCP_V_ER !�:!'O�Ko$EXTLOGo_REQ�V��I��cSIZ�o�dST�K�iU��bT�OL  �DzމR�A �d_BWD``5p�Faq�2Js�DIOq P%�es�4�f{ST�EPw��0�pOP�_DO�1FAC�TORY_TUN��Wd�yDR_GR�P 1Q�9�Ad �	{o9��0*��*�u���RH�B ��2 ���� �e9 ���m�*����z����� ׏����
��U��@�y�d�A8��?���?��?�/Ơ��
 C�0������8zc��j����3��B� � Q�A��@�33�]��33�@UU�Ty�@[�����7>�u.�>*��<���Ǒ�E�� �F@ ɢ�5W�ե��J��NJk��I'PKHu���IP�sF!{����?�  ����9�<9���896C'�6<,5�����  �H�a���{����A� ��R�ZO/�BKFEATURE� R%ap�1�ArcToo�l ���En�glish Di�ctionary���4D Stan�dard��Analog I/O���Aɰe Shif�t�rc EQ �Program �Select1�S?oftpar&�1��Weld>�ced�ures/ɯ�Co�re`Ϯ�Rampwing�utoW��wa��Updat�e��matic ?Backup�����ground E�dit����Cam�era�F
�Ce�ll��nrRn�dIm��&�omm�on calibg UI!�e�sh5��]ߋ�c�ĝ�Y�ne,����ty�sH�c��n�p�Monit�or��ntr��e�liab���DH�CP��&�ata ?Acquis��%�?iagnos����?�ocument? Viewe�'��ua��heck ?Safetyx����han|� RobF�rv�q��yս����s��FC�����x�t weav��c�h��xt. DI�O��nfi���e�nd��Err�L(t�A���s@�r�0�� Pp��FCTN �Menu�����T�P In��fac\����Gen�lsÏEq Lv����p� Mask Ex5c��g�HT��?��xy Sv��i�gh-Spe��S�kiX�m���mmounic��on��Hour����:��^��conn��2r�ncr��stru�Ҳ��KAREL �Cmd. L��u�a�Run-Ti�Env�����u+��s��S/W��License�����W�Book(S�ystem)��M�ACROs,2/�Offse��MM�R���s�Mech/Stop>�tJ�Y�"9iR�"ˍx�������od �wit�����h�.���O�ptm�a?�fi�l��`gh9ul�ti-T��ƿ�P?CM fun�i)�oV��ĉ-Regei.r��l&ri��1Fy+�&�NuE�Y�<�(C�AdjuF �.xC�#�=tatu�!�-?����RDM��o}tϰscoveر&i5em�4�n�i5pu2��	��uesL��7o�����SNPgX b���SN���Cli���>#���r�׳O� ����5ozt��ssag�� �5.���?�` ��Q�zN/I���EMIL�IB�O�BP Fi�rm�NP��Acyc�
�TPTX4��DelnQ�O�A���M�Mor�0 Si�mula��EVu��P��|J�!��&�>�ev.�E��ri���_USB pYo^�p�iPK�a����Unexcept����0�$�U����VC"t�rQH�VU�6b��OGeKAkS�0SC\UyoSUI��W�<b(�lb PlD6�n ��h�d ���w�t��|6 u�V�oCwGr{idy1play=}(�@��WwR-b.�9�-10iA/7L�MAlarm �Cause/�0e}dٸAscii>��Load���zUp�l�p��l˰��Gu���/�P���yc���� �P����RA��PC��i���`��l�p83c��NRT�z���Online HelX�m&��l&� �!��qtr��64MB� DRAM���F�RO(�Z�t� .���mai��KŅL�Sup�R*!�)��K���croE<t3E��tAfrt��t3��� <������=�4�F�s� j�|�������̯֯� ���9�0�B�o�f�x� ������ȿҿ����� 5�,�>�k�b�tϡϘ� �����������1�(� :�g�^�pߝߔߦ��� ������ �-�$�6�c� Z�l��������� ����)� �2�_�V�h� ���������������� %.[Rd�� ������! *WN`���� ����//&/S/ J/\/�/�/�/�/�/�/ �/�/??"?O?F?X? �?|?�?�?�?�?�?�? OOOKOBOTO�OxO �O�O�O�O�O�O__ _G_>_P_}_t_�_�_ �_�_�_�_oooCo :oLoyopo�o�o�o�o �o�o	 ?6H ul~����� ���;�2�D�q�h� z�����ˏԏ��� 
�7�.�@�m�d�v��� ��ǟ��П�����3� *�<�i�`�r�����ï ��̯����/�&�8� e�\�n���������ȿ �����+�"�4�a�X� jτώϻϲ������� ��'��0�]�T�f߀� �߷߮���������#� �,�Y�P�b�|��� �����������(� U�L�^�x��������� ������$QH Zt~����� � MDVp z������/ 
//I/@/R/l/v/�/ �/�/�/�/�/??? E?<?N?h?r?�?�?�? �?�?�?OOOAO8O JOdOnO�O�O�O�O�O �O_�O_=_4_F_`_ j_�_�_�_�_�_�_o �_o9o0oBo\ofo�o �o�o�o�o�o�o�o 5,>Xb��� ������1�(� :�T�^����������� ʏ��� �-�$�6�P� Z���~�������Ɵ� ���)� �2�L�V��� z�������¯���� %��.�H�R��v��� ����������!�� *�D�N�{�rτϱϨ� ����������&�@� J�w�n߀߭ߤ߶��� ������"�<�F�s� j�|���������� ���8�B�o�f�x� ������������ 4>kbt�� ����0 :g^p���� ��	/ //,/6/c/ Z/l/�/�/�/�/�/�/ ?�/?(?2?_?V?h?��?    �H541�3�12޳6R782�750޴5J614�776^�5AWSP�71�7�RCR�88�6TU��6J545�8�6V�CAM�5CLIOvPFRIOGUIF�6=66GCMSC�H�6�STYL�72FC�NRE�652�6R�63�7SCH�5DwOCV�FCSU�5�ORSFR869��70�788�6EI�O�FR54�6R6=9�6ESET,GG�JIWMG�5MA{SK�5PRXY�HM7�6OC[F`P3,H��6`P�8�853VH��XLCH�VOPLn{VJ50�VPS
gcMC�7`cW55�6�MDSWHg�WOP�WMPR[F�@�VP.�6PCMsG0�g`P��750�g517G5u1�h07FPRSWW�69�VFRDOFR�MCN�FXH93��6SNBAtG�WSHLB�FMNw�@�G�NN�X2�6HTC��6TMI�F�0VT{PA�FTPTX�v#ELv`W8�7�0�6J95FTUTv�W95�VUEC�VwUFROFVCC'��OFVIP�FCS�C�v�@Ih�6WE]B�6HTT�76�G�WIOc�CG��I�Gb�IPGS��R�C�FH77�766�7FR7JWR�hR5U3�88�h2�VR�Y�64W54��66��6|@�6NVDWVDu0R�Fu�CTO+G�NN�VOL�HENuD�6L2�FVR�E �8ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� ����������
��.� @�R�d�v����� ��������*�<�N� `�r������������� ��&8J\n �������� "4FXj|� ������// 0/B/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�? �?�?OO(O:OLO^O pO�O�O�O�O�O�O�O  __$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv���� �����*�<�N� `�r���������̏ޏ ����&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��� ����į֯������0�B�T�f�x������  H54�1����2��R78�2��50��J61�4�76��AWSuPȻ1�RCR���8�TU�J54y5��VCAM��oCLIO��RI���UIFȺ6f�CM�SC���STYLz�2G�CNREȺ�52�R63ǻS{CH��DOCVH�wCSU��ORS7ʯR869�0��8�8��EIO��R5�4׺R69�ES�ETX�&�J%�WM�G��MASK��P�RXY��7��OC����3X�׺�����53��H��LCH�'�OPL�J506g�PS��MC������55��MDSW�(�V�OPV�MPR���4�G���PCMb��0������50w�[51g�51��0gʷPRS��69G�F{RD��RMCN���u�H93�SNByA�ˆ�SHLB�ʱM�4�'�NN��2��HTC�TMI���԰��TPA��T7PTX�
EL7
����8ֻ԰��J95nG�TUTW�95G�wUEC'�UFR���VCC�O7�VI�P��CSCe�I�����WEB�HTuT�6&�WIO��CG&+IG�IP�GSX*RC��H7m7ǻ66g�R7��]R��R53��8���2g�R��64��5�4�+66������N[VD��D06;Fe<�CTOW�NNG�O]L��ENDȺL�FVR�ɗ��?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ�������� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o o&o8oJo\ono�o�o �o�o�o�o�o�o" 4FXj|��� ������0�B� T�f�x���������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� ���$�6�H�Z�l�~������STD��LANG����Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O�as�����R{BT��OPTN���,>PbDPN��z���� �����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&?�8?J?\?n?�?�:9�9�5�$FEAT�_ADD ?	�����1�0  	�8�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ��������� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� ����������&�8� J�\�n����������4DEMO R�9?   �8�� ��2);h_q ������� .%7d[m�� ������*/!/ 3/`/W/i/�/�/�/�/ �/�/�/�/&??/?\? S?e?�?�?�?�?�?�? �?�?"OO+OXOOOaO �O�O�O�O�O�O�O�O __'_T_K_]_�_�_ �_�_�_�_�_�_oo #oPoGoYo�o}o�o�o �o�o�o�oL CU�y���� ���	��H�?�Q� ~�u�������؏Ϗ� ���D�;�M�z�q� ������ԟ˟ݟ
�� �@�7�I�v�m���� ��Яǯٯ����<� 3�E�r�i�{�����̿ ÿտ����8�/�A� n�e�wϑϛ��Ͽ��� �����4�+�=�j�a� sߍߗ��߻������� �0�'�9�f�]�o�� �������������,� #�5�b�Y�k������� ����������(1 ^Ug����� ���$-ZQ c}������ � //)/V/M/_/y/ �/�/�/�/�/�/�/? ?%?R?I?[?u??�? �?�?�?�?�?OO!O NOEOWOqO{O�O�O�O �O�O�O___J_A_ S_m_w_�_�_�_�_�_ �_oooFo=oOoio so�o�o�o�o�o�o B9Keo� �������� >�5�G�a�k������� Ώŏ׏����:�1� C�]�g�������ʟ�� ӟ ���	�6�-�?�Y� c�������Ư��ϯ�� ��2�)�;�U�_��� ����¿��˿���� .�%�7�Q�[ψ�ϑ� �ϵ���������*�!� 3�M�W߄�{ߍߺ߱� ��������&��/�I� S��w������� ����"��+�E�O�|� s��������������� 'AKxo� ������ #=Gtk}�� ����///9/ C/p/g/y/�/�/�/�/ �/�/?	??5???l? c?u?�?�?�?�?�?�? OOO1O;OhO_OqO �O�O�O�O�O�O
__ _-_7_d_[_m_�_�_ �_�_�_�_o�_o)o 3o`oWoio�o�o�o�o �o�o�o%/\ Se������ ���!�+�X�O�a� ������ď��͏��� ��'�T�K�]����� ������ɟ������ #�P�G�Y���}����� ��ů������L� C�U���y��������� ������H�?�Q� ~�uχϴϫϽ����� ����D�;�M�z�q� �߰ߧ߹�������	� �@�7�I�v�m��� �����������<� 3�E�r�i�{������� ������8/A new����� ��4+=ja s������� /0/'/9/f/]/o/�/ �/�/�/�/�/�/�/,? #?5?b?Y?k?�?�?�? �?�?�?�?�?(OO1O ^OUOgO�O�O�O�O�O �O�O�O$__-_Z_Q_ c_�_�_�_�_�_�_�_ �_ oo)oVoMo_o�o �o�o�o�o�o�o�o %RI[������}   �x�	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i�{�������ÿ տ�����/�A�S� e�wωϛϭϿ����� ����+�=�O�a�s� �ߗߩ߻�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C Ugy����� ��	-?Qc u������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s��������������  ������ 1CUgy��� ����	-? Qcu����� ��//)/;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?m?? �?�?�?�?�?�?�?O !O3OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_e_w_�_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹������� ��%�7�I�[�m�� ������������� !�3�E�W�i�{�����P������������ ��#5GYk} ������� 1CUgy�� �����	//-/ ?/Q/c/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{�������y�$F�EAT_DEMO�IN  �t�����p�tIND�EX����pI�LECOMP �S���M����uC�SETU�P2 TM�~W��  N ���@�_AP2BCK� 1UM�  #�)�x��ŋ%����pP�׏��u��@� Ϗd��q���)���M� ��������<�N�ݟ r������7�̯[�� ���&���J�ٯn��� ���3�ȿڿi����� "�4�ÿX��|�ω� ��A���e���ߛ�0� ��T�f��ϊ�߮��� O���s����>��� b��߆��'��K��� ������:�L���p� ���#�����Y���}� $��H��l~ �1��g��  �-V�z	�� ?�c�
/�./� R/d/��//�/;/�/��/\���P�� 2>��*.VR�/3?� *6?\?�#b?�?�p%0PC�?�?� OFR6:�?�>r?O�;T+�+O=O�5(O�gL��?�Oo&*.F ?�O�!	�3�O�LqzO_�KSTM_ D_�2�00_o]�O�_�KH`_�_UW�_q_�_o�JGIF"oLoWU�8o�_o�o�JJPG �o�oWU�oyo�o �:#JS*S� �cA��o%
JavaS�cript�oC�Sp�VV�� %�Cascadi�ng Style Sheets��u 
ARGNAMOE.DT2��,ZP�\F��fqv���3�>v�DISP*}�`��ZPʏ
��������
�TPEINS.X3ML:��:\N���n�Custom Toolbar�����PASSWOR�D��.FRS:�\ҟ�� %Pa�ssword Config�n/\� �U����/��E�گ� {����4�F�կj��� ���/�ĿS��w�� ϭ�B�ѿf�x�Ϝ� +�����a��υ�ߩ� ��P���t��mߪ�9� ��]�����(��L� ^��߂���5�G��� k� �����6���Z��� ~������C�����y� ��2����h��� ��Q�u
 �@�dv�) �M_��/�/ N/�r//�/�/7/�/ [/�/?�/&?�/J?�/ �/�??�?3?�?�?i? �?�?"O4O�?XO�?|O �OO�OAO�OeOwO_ �O0_�O)_f_�O�__ �_�_O_�_s_oo�_ >o�_bo�_o�o'o�o Ko�o�o�o�o:L �op�o��5�Y �}�$��H��A� ~����1�Ə؏g��� �� �2���V��z�	� ���?�ԟc�͟
��� .���R�d�󟈯��� ��M��q������<� ˯`��Y���%���I� ޿��ϣ�8�J�ٿ�n�����!�3��ϫ���$FILE_DG�BCK 1U�������� < �)
S�UMMARY.DyG��~�MD:��F���Diag� Summary�G�T�
CONSLOG<��1ъ���Y��Console� log��S�	T�PACCN��%�%��J�U�TP A�ccountin���T�FR6:I�PKDMP.ZI	P~��
����V�f��Exceptio�n���2�MEMCHECK@��5�V����Memory� DataW����/YF)	FTP��߮�=���a���m�ment TBD�����L =�)�ETHERNET���|��^Y�E�thernet ~��figura���Z���DCSVRF��������g�%��  verify� all���M{+��DIFF�p��eh�%�diffg� CHG01\CU`��}/*f�2���n/y/!/¯3d/K/]/�/ ��/?�&VTR�NDIAG.LS�?�/�/v?i�61 ~^�nosticw?���T6a)UPDATES.�0��?�FRS:\��?�=Z�Upda�tes List��?|�PSRBWLOD.CM*O~��2�>O�?��PS_RO�BOWEL��R�>b1HADOWl?Q?�c? _g�Shad�ow Changses_��q�BNOTI��O�O�_�e�Notifi�c�'_��+@AG `��_���_��
o3oZ� Wo�_{o�oo�o@o�o �ovo�o/A�oe �o���N�r ���=��a�s�� ��&���͏\�񏀏� ��"�K�ڏo������� 4�ɟX������#��� G�Y��}����0��� ׯf������1���U� �y������>�ӿ� t�	Ϙ�-ϼ�:�c�� ��ϫϽ�L���p�� ߦ�;���_�q� ߕ� $߹�H�����~��� 7�I���m��ߑ��2� ��V������!���E� ��R�{�
���.����� d�����/��S�� w��<�`� �+�Oa�� ��J�n// �9/�]/�j/�/"/ �/F/�/�/|/?�/5? G?�/k?�/�?�?0?�? T?�?x?�?O�?CO�? gOyOO�O,O�O�ObO �O�O_-_�OQ_�Ou_ _�_�_:_�_^_�_o �_)o�_Mo_o�_�oo �o�oHo�olo�o 7�o[�o� � D��z��3�E� �i�������ÏR� �v�����A�Џe� w����*���џ`��� �����&�O�ޟs�� ����8�ͯ\����� '���K�]�쯁�����4���ۿ���$FI�LE_FRSPRT  ��Ű�����MDONLY 1�UŽ� 
 ��)MD:_V�DAEXTP.Z�ZZ⿓�j�y��6%NO Ba�ck file <DϽ�S�6p��� Z��ϸ���%�j�I��� m��ߣ�2�����h� �ߌ�!�3���W���{� 
���@���d���� ��/���S�e����� ����N���r��� =��a����&� J����9K~��VISBCK"�|�1�*.VDL|�FR:\e�ION\DATA�\�'Vision VD�� ��
//2@/*d/ �u/�/)/�/M/�/�/ �/?�/<?�/�/r?? �?�?c?�?[?�??O &O�?JO�?nO�OO�O 3O�OWOiO�O�O"_4_ �OX_�O|__�_�_A_ �_e_�_o�_0o�_To��_�_�o�LUI_�CONFIG �V�x�k '$ sc'�{��o��o"4FTy�`|x|o~�����| l���/�A��R� w���������V���� ��+�=�ԏa�s��� ������R�ߟ��� '�9�П]�o������� ��N�ۯ����#�5� ̯Y�k�}�������J� ׿�����1�ȿU� g�yϋϝ�4Ϯ����� ��	�߲�?�Q�c�u� �ߙ�0߽�������� ��;�M�_�q��� ,������������ 7�I�[�m����(��� ����������3E Wi{�$��� ���
/ASe w������ �/+/=/O/a/s/
/ �/�/�/�/�/�/�/? '?9?K?]?o??�?�? �?�?�?�?�?O#O5O GOYOkOO�O�O�O�O �O�O�O__1_C_U_ �Of_�_�_�_�_�_j_ �_	oo-o?oQo�_uo �o�o�o�o�ofo�o );M�oq�� ���b���%� 7�I��m�������� ǏZ�����!�3�E��Ոa�|�$FL�UI_DATA �W���v��فh�RESULT 2Xv���� �T��/wizard�/guided/�steps/ExpertQ�֟��� ��0�B�T�f�x�������Conti�nue with{ G��ance�� ӯ���	��-�?�Q��c�u����� _�-�`�v���0 �`း�x�w�ع���ps��#�5�G�Y�k� }Ϗϡϳ������Ϩ� ��"�4�F�X�j�|� �ߠ߲���������ؿ�ʿܿ���torch�p����� ������ ��$�6��� Z�l�~����������� ���� 2D���_9�K�wproc _�����0 BTfx�I��� ���//,/>/P/ b/t/�/�/Wi�/��������Time?US/DST�/*? <?N?`?r?�?�?�?�?��?�?��Disabl��O%O7OIO[O mOO�O�O�O�O�O�N_�ـ�/�/�/�/�/224?z_�_ �_�_�_�_�_�_
oo .o�?�?dovo�o�o�o �o�o�o�o*<��O__1_󷩟��Region?�� ���(�:�L�^�p������America���Ώ���� �(�:�L�^�p�����Jqy��j̟��
2EdiZ���"�4�F� X�j�|�������į֯�� Touch �Panel � �(recommen	�)�)�;�M�_� q���������˿ݿ�������� ����
2acces��uχϙ� �Ͻ���������)���Connec�t to Network8�o߁ߓ� �߷����������#�5�X�t�6���!J�0Introduct������� ��'�9�K�]�o��� ��������������#5GYk}� �/b���HR�� &8J\n�� �������/"/ 4/F/X/j/|/�/�/�/��/�/Fx� ��
���~ ?*?�Q? c?u?�?�?�?�?�?�? �?OO)O�MO_OqO �O�O�O�O�O�O�O_ _%_�/�/??|_>? �_�_�_�_�_�_o!o 3oEoWoio{o:O�o�o �o�o�o�o/A Sew�H_Z_l_� �_���+�=�O�a� s���������͏�o� ��'�9�K�]�o��� ������ɟ۟���  ��G�Y�k�}����� ��ůׯ�����ޏ 0�U�g�y��������� ӿ���	��-��N� �r�4��ϫϽ����� ����)�;�M�_�q� �ߔϧ߹�������� �%�7�I�[�m��>� ��b���������!� 3�E�W�i�{������� ��������/A Sew����� ��������Oa s������� //'/��K/]/o/�/ �/�/�/�/�/�/�/? #?�D?h?z?>/�? �?�?�?�?�?OO1O COUOgOyO8/�O�O�O �O�O�O	__-_?_Q_ c_u_4?~?X?�_�_�? �_oo)o;oMo_oqo �o�o�o�o�o�O�o %7I[m� ����_�_�_�� �_E�W�i�{������� ÏՏ������oA� S�e�w���������џ ��������� p�2�������ͯ߯� ��'�9�K�]�o�.� ������ɿۿ���� #�5�G�Y�k�}�<�N� `��τ�������1� C�U�g�yߋߝ߯��� ������	��-�?�Q� c�u�������� �ϲ����;�M�_�q� �������������� ��$I[m� ������! ��B�f(���� ����////A/ S/e/w/��/�/�/�/ �/�/??+?=?O?a? s?2�?V�?z�?�? OO'O9OKO]OoO�O �O�O�O�O�/�O�O_ #_5_G_Y_k_}_�_�_ �_�_�?�_�?
o�?�_ CoUogoyo�o�o�o�o �o�o�o	�O?Q cu������ ����_8��_\�n� 2������ˏݏ�� �%�7�I�[�m�,�� ����ǟٟ����!� 3�E�W�i�(�r�L��� ���������/�A� S�e�w���������~� �����+�=�O�a� sυϗϩϻ�z�į�� ���ԯ9�K�]�o߁� �ߥ߷���������� п5�G�Y�k�}��� ��������������� ���d�&ߋ������� ������	-?Q c"������ �);M_q 0�B�T��x���/ /%/7/I/[/m//�/ �/�/t�/�/�/?!? 3?E?W?i?{?�?�?�? �?���O�/OAO SOeOwO�O�O�O�O�O �O�O_�/_=_O_a_ s_�_�_�_�_�_�_�_ oo�?6o�?ZoO�o �o�o�o�o�o�o�o #5GYk|o�� �������1� C�U�g�&o��Jo��no ӏ���	��-�?�Q� c�u���������|� ���)�;�M�_�q� ��������x�گ���� ��¯7�I�[�m���� ����ǿٿ����Ο 3�E�W�i�{ύϟϱ� ���������ʯ,�� P�b�&ωߛ߭߿��� ������+�=�O�a�  υ���������� ��'�9�K�]��f� @ߊ���v������� #5GYk}�� �r����1 CUgy���n� �����/��-/?/Q/ c/u/�/�/�/�/�/�/ �/?�)?;?M?_?q? �?�?�?�?�?�?�?O ����XO/O�O �O�O�O�O�O�O_!_ 3_E_W_?{_�_�_�_ �_�_�_�_oo/oAo Soeo$O6OHO�olO�o �o�o+=Oa s���h_��� ��'�9�K�]�o��� ������vo�o�o���o #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	�ȏ*��N� �u���������Ͽ� ���)�;�M�_�p� �ϕϧϹ�������� �%�7�I�[��|�>� ��b����������!� 3�E�W�i�{���� p���������/�A� S�e�w�������l��� �����߶�+=Oa s������� ��'9K]o� ���������  /��D/V/}/�/�/ �/�/�/�/�/??1? C?U?y?�?�?�?�? �?�?�?	OO-O?OQO /Z/4/~O�Oj/�O�O �O__)_;_M___q_ �_�_�_f?�_�_�_o o%o7oIo[omoo�o �obO�O�O�o�o�O! 3EWi{��� �����_�/�A� S�e�w���������я ����o�o�o�oL� s���������͟ߟ� ��'�9�K�
�o��� ������ɯۯ���� #�5�G�Y��*�<��� `�ſ׿�����1� C�U�g�yϋϝ�\��� ������	��-�?�Q� c�u߇ߙ߫�j�|��� �߲��)�;�M�_�q� ������������  �%�7�I�[�m���� �������������� ��B�i{��� ����/A Sdw����� ��//+/=/O/ p/2�/V�/�/�/�/ ??'?9?K?]?o?�? �?�?d�?�?�?�?O #O5OGOYOkO}O�O�O `/�O�/�O�/�O_1_ C_U_g_y_�_�_�_�_ �_�_�_�?o-o?oQo couo�o�o�o�o�o�o �o�O�O8Joq �������� �%�7�I�om���� ����Ǐُ����!� 3�E�N(r���^ ß՟�����/�A� S�e�w�����Z���ѯ �����+�=�O�a� s�����V���z�Ŀ� ���'�9�K�]�oρ� �ϥϷ������Ϭ�� #�5�G�Y�k�}ߏߡ� �������ߨ���̿޿ @��g�y������ ������	��-�?��� c�u������������� ��);M�� 0�T���� %7I[m� P������/!/ 3/E/W/i/{/�/�/^ p��/�??/?A? S?e?w?�?�?�?�?�? �?��?O+O=OOOaO sO�O�O�O�O�O�O�O �/_�/6_�/]_o_�_ �_�_�_�_�_�_�_o #o5oGoX_ko}o�o�o �o�o�o�o�o1 C_d&_�J_�� ���	��-�?�Q� c�u�����Xo��Ϗ� ���)�;�M�_�q� ����T��xڟ��� �%�7�I�[�m���� ����ǯٯ믪��!� 3�E�W�i�{������� ÿտ翦��ʟ,�>� �e�wωϛϭϿ��� ������+�=���a� s߅ߗߩ߻������� ��'�9���B��f� ��RϷ���������� #�5�G�Y�k�}���N� ����������1 CUgy�J��n� ����	-?Q cu������ ��//)/;/M/_/q/ �/�/�/�/�/�/�� ��4?�[?m??�? �?�?�?�?�?�?O!O 3O�WOiO{O�O�O�O �O�O�O�O__/_A_  ??$?�_H?�_�_�_ �_�_oo+o=oOoao so�oDO�o�o�o�o�o '9K]o� �R_d_v_��_�� #�5�G�Y�k�}����� ��ŏ׏�o���1� C�U�g�y��������� ӟ埤��*��Q� c�u���������ϯ� ���)�;�L�_�q� ��������˿ݿ�� �%�7���X��|�>� �ϵ����������!� 3�E�W�i�{ߍ�L��� ����������/�A� S�e�w��HϪ�l��� �ϒ���+�=�O�a� s��������������� '9K]o� ����������  2��Yk}�� �����//1/ ��U/g/y/�/�/�/�/ �/�/�/	??-?�6 Z?�?F�?�?�?�? �?OO)O;OMO_OqO �OB/�O�O�O�O�O_ _%_7_I_[_m__>? �?b?�_�_�?�_o!o 3oEoWoio{o�o�o�o �o�o�O�o/A Sew����� �_�_�_�_(��_O�a� s���������͏ߏ� ��'��oK�]�o��� ������ɟ۟���� #�5����z�<��� ��ůׯ�����1� C�U�g�y�8������� ӿ���	��-�?�Q� c�uχ�F�X�j��ώ� ����)�;�M�_�q� �ߕߧ߹��ߊ���� �%�7�I�[�m��� ������������ ��E�W�i�{������� ��������/@� Sew����� ��+��L� p2������� //'/9/K/]/o/�/ @�/�/�/�/�/�/? #?5?G?Y?k?}?<�? `�?��?�?OO1O COUOgOyO�O�O�O�O �O�/�O	__-_?_Q_ c_u_�_�_�_�_�_�? �_�?o&o�OMo_oqo �o�o�o�o�o�o�o %�OI[m� �������!� �_*ooN�x�:o���� ÏՏ�����/�A� S�e�w�6������џ �����+�=�O�a� s�2�|�V���ʯ��� ��'�9�K�]�o��� ������ɿ������ #�5�G�Y�k�}Ϗϡ� ���τ��������ޯ C�U�g�yߋߝ߯��� ������	��ڿ?�Q� c�u��������� ����)������n� 0ߕ����������� %7I[m,� ������! 3EWi{:�L�^� �����////A/ S/e/w/�/�/�/�/~ �/�/??+?=?O?a? s?�?�?�?�?�?��? �O�9OKO]OoO�O �O�O�O�O�O�O�O_ #_4OG_Y_k_}_�_�_ �_�_�_�_�_oo�? @oOdo&O�o�o�o�o �o�o�o	-?Q cu4_����� ���)�;�M�_�q� 0o��To��xoz��� �%�7�I�[�m���� ����ǟ�����!� 3�E�W�i�{������� ï��䯦���ޟA� S�e�w���������ѿ �����؟=�O�a� sυϗϩϻ������� ��ԯ���B�l�.� �ߥ߷���������� #�5�G�Y�k�*Ϗ�� ������������1� C�U�g�&�p�Jߔ��� ������	-?Q cu����|�� �);M_q ����x������� /��7/I/[/m//�/ �/�/�/�/�/�/?� 3?E?W?i?{?�?�?�? �?�?�?�?OO��  /bO$/�O�O�O�O�O �O�O__+_=_O_a_  ?�_�_�_�_�_�_�_ oo'o9oKo]ooo.O @ORO�ovO�o�o�o #5GYk}�� �r_�����1� C�U�g�y��������� �o⏤o��o-�?�Q� c�u���������ϟ� ���(�;�M�_�q� ��������˯ݯ�� �ҏ4���X����� ����ǿٿ����!� 3�E�W�i�(��ϟϱ� ����������/�A� S�e�$���H���l�n� ������+�=�O�a� s�����z����� ��'�9�K�]�o��� ������v������� ��5GYk}�� �������1 CUgy���� ���	/����6/ `/"�/�/�/�/�/�/ �/??)?;?M?_? �?�?�?�?�?�?�?O O%O7OIO[O/d/>/ �O�Ot/�O�O�O_!_ 3_E_W_i_{_�_�_�_ p?�_�_�_oo/oAo Soeowo�o�o�olO~O �O�O�O+=Oa s������� ��_'�9�K�]�o��� ������ɏۏ���� �o�o�oV�}����� ��şן�����1� C�U��y��������� ӯ���	��-�?�Q� c�"�4�F���j�Ͽ� ���)�;�M�_�q� �ϕϧ�f�������� �%�7�I�[�m�ߑ� �ߵ�t��ߘ��߼�!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ������(��L� s������� '9K]�� �������/ #/5/G/Y/z/<�/ `b/�/�/�/??1? C?U?g?y?�?�?�?n �?�?�?	OO-O?OQO cOuO�O�O�Oj/�O�/ �O_�?)_;_M___q_ �_�_�_�_�_�_�_o �?%o7oIo[omoo�o �o�o�o�o�o�o�O_ �O*T_{��� ������/�A� S�ow���������я �����+�=�O� X2|���h͟ߟ� ��'�9�K�]�o��� ����d�ɯۯ���� #�5�G�Y�k�}����� `�r����������1� C�U�g�yϋϝϯ��� �����϶��-�?�Q� c�u߇ߙ߽߫����� ���Ŀֿ�J��q� ������������ �%�7�I��m���� ������������! 3EW�(�:�^� ����/A Sew��Z��� ��//+/=/O/a/ s/�/�/�/h�/��/ �?'?9?K?]?o?�? �?�?�?�?�?�?�?? #O5OGOYOkO}O�O�O �O�O�O�O�O�/_�/ @_?g_y_�_�_�_�_ �_�_�_	oo-o?oQo Ouo�o�o�o�o�o�o �o);M_n 0_�T_V���� �%�7�I�[�m���� ��boǏُ����!� 3�E�W�i�{�����^ ���������/�A� S�e�w���������ѯ ������+�=�O�a� s���������Ϳ߿� ����ԟ�H�
�oρ� �ϥϷ���������� #�5�G��k�}ߏߡ� ������������1� C��L�&�p��\��� ������	��-�?�Q� c�u�����X߽����� ��);M_q ��T�f�x����� %7I[m� �������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/���>?  e?w?�?�?�?�?�? �?�?OO+O=O�aO sO�O�O�O�O�O�O�O __'_9_K_
??.? �_R?�_�_�_�_�_o #o5oGoYoko}o�oNO �o�o�o�o�o1 CUgy��\_� �_��_	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�q� ��������˟ݟ ��4��[�m���� ����ǯٯ����!� 3�E��i�{������� ÿտ�����/�A�  �b�$���H�JϿ��� ������+�=�O�a� s߅ߗ�V��������� ��'�9�K�]�o�� ��Rϴ�v������� #�5�G�Y�k�}����� ����������1 CUgy���� ��������<�� cu������ �//)/;/��_/q/ �/�/�/�/�/�/�/? ?%?7?�@d?�?��1�$FMR2_�GRP 1Y�5�� ��C4  B�N 	� N �?�<�0E�� F@ �2ǂ5WEF:�0J���NJk�I'�PKHu��IP��sF!��M?ǀ  JOF<�09��<9�8�96C'6<�,5��MAg�  �O�KBH�3�B��0�@�A@�3]3�B�33F<�4x�O]�0@UUTZ�@�@+PMJ)>u.��>*��<����M=[�B=����=|	<��K�<�q�=��mbN��8��x	7H<8��^6�Hc7��x2_�__�_�_�_�o o9oL'�2_CF�G Z�;T �Do�o�o�oKkNO� �:
F0��a �`JlRM_C�HKTYP  ��1N �0�0u0�1RO=M�`_MIN pN#W��,p��@X�0�SSB[c[�5 �6YN%�Psy�QeTP_D�EF_O@N$|�3�wIRCOM�`���$GENOV_RD_DO!vW!n�}THR!v d�u�d�t_ENB� ��pRAVC�3\�BwMp ��5F�s  G!� G�Ƀ�I�C�I(i J���ohu��N"�0"p�ÅF���F �VD�OU�0b�<�aq�8�r�5<)p ^M6���.�P�~�~N#C�  D��`�ȟ؜^HŖB��1�Œ�9!��E�SMT®3cR��0Op���$�HOSTC[b1d��9Np�W/�0 3MC���y�L&  27.0ɠ=1��  e���� ��,�:��]�o���𓿶�M�G�	anonymoul�ؿ꿀��� �2�x��0E� E˧�����ݯ������ ���I�&�8�J�\�� �ǿ�߶�������3� ��W�i�F�}ߟ�]�� ������������ 0�S�ߛ�x������� ����+�=�?�,s� Pbt����� ��']�L^ p���������  /G$/6/H/Z/�~/ �/�/�/�/�k/1?  ?2?D?V?���� �/�?	/�?�?
OO.O u/ROdOvO�O�O�?�/ ?�O�O__*_q?�? �?r_�O�_�?�_�_�_ �_�O�_&o8oJo\o_ �o�O�o�o�o�o�o3_ E_W_i_ko=�_|� ���o���� 0�S�o�ox����������-�[�ENT 1=e� P!I��  *���2�!� V��z�=���a����� ӟ�����ߟ@��d� '���K�]�����⯥� �ɯ*����`�#��� G���k�̿��ſ�� &��J��n�1�z�U� ���ϋ��ϯ����4� ��X��-ߎ�Q߲�u���ߙ�QUICCA0�߿���2���13��!����2��_�q����!ROUTE�R�����"�!P�CJOG#���!�192.168�.0.10����C�AMPRTs�O�!�c�1l����RT������ׄNAM�E !�!R�OBO��S_C�FG 1d� ��Aut�o-starte�dtFTP% �<>��r� /A�ew��� �R��//+/�#�v����/� ��/�/�/�/?�&? 8?J?\?n?�/?�?�? �?�?�?�?'9 }?jO�/�O�O�O�O�O �?�O__0_B_eO�O x_�_�_�_�_�_O+O =OoQ_>o�Oboto�o �o__�o�o�o�o'o �o#L^p���_ �_�_o �Go$�6� H�Z�l�3������Ə ؏�}�� �2�D�V� h�������ԟ� ��
��.����d�v� ��������Q����� �*�q���������{� ݟ��̿޿��ɯ&� 8�J�\�nϑ�Ϥ϶� ��������E�W�i�� }�j߱��ߠ߲����� ������0�S�T��߀x������T( _?ERR f2
�����PDUSIZ � b�^�����>�WRD ?�qB��  ?guest`�P��b�t�������!SC�DMNGRP 2�gq����B�b�[$`�K�� �	P01.02� 8'�   ���  �� @  
=� ����wG�*����uG �����7��k����4�w ���B(Ї7�)������ r�������y��-�"BC�l�
d�-?Q��_GROUU��h�������	���QUPD'  >������TYf ����T�TP_AUTH �1i�� <!iPendan���,.k�!K?AREL:*,/5/G-KC\/l/~/T �VISION �SET��/�/b� R"�/�/?Q#/??G? A?�?e?w?�?�?�>�CTRL j�����Eb�
b�F�FF9E3�?@��FRS:DEFA�ULT:LFA�NUC Web ?Server:J(B �8�J��<�O�O�O�O��O_��WR_CONFIG k��� :O��IDL_CPU_PCY@�b�B�C�xP BH^UMINi\(�|U?GNR_IO����b���`PNPT_S_IM_DO�V�[�STAL_SCR�N�V ��INT�PMODNTOL8�W�[�ARTY�XxQ�V� �EN� �U��\TOLNK 1l��L��o�o�o�o��o�o�odbMAST�E�P�dbSLAV�E m��uRA?MCACHE
b}O!O_CFGL�ccdsUO�o`rC�YCLK~uS@_A�SG 1n��*�
 �o���'�9� K�]�o���������ɏ�ۏ�k�rNUM����
`rIPI[wR?TRY_CNY@�R@��`r�Q��a���1 `r�piro*~D����D�`PSDT_I�SOLC  ����$J23_DeSLdN��OG��1p*{<��<zPE�?��,��?�	߂�Q�������ʯ��� ��$�`��Οؘ��PeqC�ޒP�BpECMo�UKANJI_p �_��Z ?MON q�_b�y���&�8�J�H�X"��r;\Fl�<����CL_L�P��$���EYLOGG+INlpD�������$LANGU�AGE �F;beSD ���LGjq�s�y`a �*b�xC�G�J@~P��b�'0_�b�;�b�=MH ;���
��(UT1:\ZϤߥ�߷����� ����#�L�G�Y�~��(����LN_D?ISP t*qؘ��~���OCboRD�z�S�A�OGB?OOK u'���`������Xp� i�{�������O*3�K���F	+�r١B�s�(:s����_B�UFF 1vom?�J@tD� B� CG�����! *WN`���������/��XD�CS x�{� =�����!��E�/�/�/�/4$IO 1y�{ ���#�0��/??(?<?L?^? p?�?�?�?�?�?�?�?  OO$O6OHO\OlO~Oh�O�O�%E�PTM��dB��O_!_3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeo�N�BSEVd����FTYP���O�o�o�otm��RSB���V>\�FL 2z�-j��e/ew�����TP�����b}�NGNAM锸%�0$UPS��G�IB���o�@�_L�OADPROG �%��%PLA�CE_SALID�A���MAXUALRM��A���F�'_PRB�f� �����C��{'����x����P 2|��W ؄	�a�
*eЃ��X��� o�����c(���ԟ� ��C�.�g�R����� �������ȯگ�� ?�*�c�u�X������� �����޿��;�M� 0�q�\ϕ�xϊ��϶� �����%��I�4�m� P�bߣߎ��߲����� ��!��E�(�:�{�f� �������������  ��S�>�w�b����������������DBG?DEF }�u!����� _LDXD�ISA+��{�#ME�MO_AP%�E {?�{
 " �~����������ISC 1~
�y�����IS�'�_�����+_MSTR �m~�SCD 1�m��./�R/=/v/a/ �/�/�/�/�/�/�/? ?<?'?L?r?]?�?�? �?�?�?�?O�?�?8O #O\OGO�OkO�O�O�O �O�O�O�O"__F_1_ j_U_g_�_�_�_�_�_ �_o�_oBo-ofoQo �ouo�o�o�o�o�o �o,P;t_� ���������:��MJPTCF/G 1��7�����[`�MIR 1e����J�@���D@ !1��Ñc�K�؏��< ��� �?�� �����C�j���N�  �I��A�c���w���ǟ������ӟ E�+�3�=���a���� ϯ��ׯ����K� ]�����f�p���̿ j�Ŀֿ����J�,� }Ϗϡ�4�V��Ϫ��� ��߮��F�,�>�`� b�p�����f�xߚ�� �����T�:�\��p� ����ߴ������ ����2�<�N�`�~��� ����������I[ ���d�v���h ����H*{ ��2T���� /�/D/*/</^/�/�n]�Kc��i� � �/[�LTARkM_�"�������"w�n�?4]�ME�TPU  ���%\�NDSP?_ADCOL25� �=>CMNTS? ~F5MST ��-��?w��!�?�4F5PO�SCFs7~>PR�PMr?�9STQ01��i�4��<#�
 AA5�AEQO_G=O_OaO sO�O�O�O�O�O�O!_ __W_9_K_�_o_�_��_�QF1SING_�CHK  V?$_MODAQ�#�i��#5v�U�5U� b�DEV 	i�	�MC:1lHSI�ZE20�-��UTA�SK %i�%$�12345678�9 �o�e�WTRI�e��i� l��% ��og�o)}���c�YPkaz�d�SE�M_INF 1���'a`)AT&FV0E02��})�qE0V1�&A3&B1&D�2&S0&C1S�0=�})ATZ���tH�)��qQ��xAY���<�����ɏۏ � ���� �Z��~�������g� ؟�������2���� h��-�?�����u�� �
�ůϟ@���d�K� ����M���q������� �˯<�s�M�r�%��� QϺ��ϳ��ϣ���&� ٿ���n߀�3Ϥ��� �߃ߍ��߹�"�	�F� X��|�/�A�S�e��� �����C�0���T���e���q����.ONIwTOR�0G ?Ek�   	EX�EC1o"��2��3���4��5���`��7*��8��9����x� \��\\\ \&\2\>\J�\V\2c2o2�{2�2�2�2��2�2�2�3�c3o3�QR_�GRP_SV 1��~{ (�Qo!�����?nt���_N���"�g�����a_DM��nn�ION_DB�`�mo!  a�� �#� w+��o  h��N �l() i-ud�1Wem//�/�!PL�_NAME !��e� �!De�fault Pe�rsonalit�y (from �FD)<"*0RR2�u 1�L68�L@P�!`
 d�??,?>?P? b?t?�?�?�?�?�?�? �?OO(O:OLO^OpO�O��2?�O�O�O�O��O__*_<_N_��< �Ox_�_�_�_�_�_�_��_oo,o>o=,��Dg_xn
go�o��P�o �o�o�o�o"4F Xj|����� �o�o��0�B�T�f� x���������ҏ��� ����P�b�t��� ������Ο������(�:�L�^�p� �Fs  GT��G�M����(������d�ͯ߮ į����u�p��H�pX�B�{�~� k� ��������οԿ�Ϡ��7�G̛�k�	�`��zόϞ�]�:�oA<)�����ϙ� A�  	٤�"�#��)2 h�?, � �� ~;� @D�  N�?�T�:�?��Vћ�A/��N�Un��;��	lf�	 �xJ���3 � �� ��< ���� ���ґK�K� ��K=*�J����J���J9�]��\������@�t�@{S�6��(EB�n������=�N��I�l�T;f�a���������* � ´  � Õ>�����T��>����ӧU�'�x`������g���j�\!�}ߑ��  {  �@* ���  ��" �F�j�d��	�'� � ���I� �  y�
Ш�:�È��?È=��;���[��( �5��n @����@���i�@�����;!P�  'f3�g�@�2��@�0@js�@w�@{�C��}C< C��\C���C��C��!!�K@���f� ��d0�B< �	�����&��Dzc�I��mX�}����( ?�� -����`�����A���0%��������?�faf!�//� W��K/]+��8��s/�*>���<�b��(���%P��(��ѮӮ�?�����x�����<�
6b<߈;�܍�<�ê<���<�^���d#?��A��U��@�|f��?fff?9��?&`0.�@�.�r2�J<?�\�~2N\����[1g� �Vն?T��?D7��5/ 
O�?.OORO=OvOaO��O�O�O�O�ȟ5F ���O_�O0_�?Q_�9�#_�_XG@ G�@0��G�� G}��s_�_�_�_�_o�o@o+oBL��Bh�AQo5o�o�m-�m �o���K_o_8�o�\n��|��b�|��#/A @|J �F���=�/ù�!A� Z���A*���x&��ߞ�?�ؽ��ď��菦��W������CP�K�CH��BZׄ���ցz�@�I�Vn(hA�� �ALffA�]��?�$�?���!�°u��æ�)�	ff���C�#�
�^���g\)�2�3�3C�
������<���G��B���L��B�s�����	�"�H����G��!G���WIYE����C�+��I�۪I�5�H�gMG�3E���RC�j=R�
��pI���G���fIV=�E<YD�S����� ۯƯد���5� �Y� D�}�h�������׿¿ ����
�C�.�@�y� dϝψ��Ϭ������� ��?�*�c�N߇�r� �ߖߨ��������)� �M�8�]��n��� �����������I� 4�m�X���|������� ������3WB {fx�������(������?�"��^�����N`��3�8��z���4Mgux�����VwQ���4p�+4�]��>/,/b/P/�/�t,�eP2P�.�a �o�/4�/??;?&;RA?H?�?l?�?�?�?  ��?�?O �?)OOMO�/�o�OnO�O�K�O�O�O�O�O __�"&_8_n_�\_�_�_�_�Z  2� Fs��GT]��V�M��B)�XV�c�J�C�pc@g� ,o��ISoeowo�o�o� �\!��WɃ�Bo�o�oz?��W�@@z�������������
 s���� �����'�9�K��]���Mq �����D��$MSK�CFMAP  ��� �VMqIq��ONR�EL  �%���CP��EXCFE�NB߇
��х��F�NC���JOGO'VLI�P�d��]d��KEY߇K�=T�_PANވf�\b���RUN;�K����SFSPDTY�� ��ӃSIGN|ߏ�T1MOT=�����_CE_G�RP 1����\>OB�6Of�x��T b���Z�ǯ~������� !�د�W��{���D� ��h�տ翞��¿� A���e�w�^ϛ�RϿ���ϸ��ϡf��QZ_�EDITܔ��уT�COM_CFG 1���XvP�b�t�}
0�_ARC_����%*�T_MN_oMODEܖ�
�UAP_CPL����NOCHECK� ?��  �%����1�C�U�g� y�������������	��ȋNO_WA�IT_Lۗ%��NMT8����O{m�o_ERR�2���CQ� �����������|� �Բ�O����|	�f����BUz��G�#��!'j³�&K2<��h?�l�%Hp����_PARAM�򙣋�	��N8��_8 =�P345?678901Rd vM������`�/%/+N7�W/�i,��/тODRD�SP��ޖ
�OFFSET_CARМ���&DIS�/�#S;_A��ARKܗ&��OPEN_FIL�E� B�v�&֎�OPTION_IO\����G0M_PRG ;%��%$*�?�>�#3WO0� ��
t �5��tN��� ����0��1	 ����1������� RG_DS�BL  ����P|LO�!RIENTkTOހ��C�Gp���a� UT_SIM_DO7��}�� �V� LCT � w�"��4v��I��S��A�_PEX���/�DR[AT�� d
��D>� UP ��N^p!��C_U_2r@SubAq�RH�W]�$��2��L68L�@P�C
 d}/�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6��2�_fx���� ����}U2�D� V�h�z�������ԏ ������"�2�pP2�X���PE��������� ʟܟ� ��$�6�H� Z�l�~���_�q�Ưد ���� �2�D�V�h� z�������¿Կ���� 
��.�@�R�d�vψ� �ϬϾ������������O'�W�i��C{$�ߙ�~߼���<�@<�|/���1����  �P�F�X�j������$�sQ����	�`:�4�F�X���:�o{Av�������%�A�  ���T�P�O)P1�[��v�T"��, �D[0�� @D�  ��:��?�D��� H;�	l�	� �xJf �9:] � �< ��| ��0�$�H(���H3k7HSM�5G�22G���GN�3�HI�X��$�Cfp@ap@B���,Q#ã0��s@�4*>*�*�9/�A�q�½{q�ª3��Pd ���%�$���;$�}��@{  @k@}�P0�  ��0��&$�"/P%	'�� � @"I� �  ���f=���d/v+����  ���n @�"�A�/'+B����9N|@?  'R0&4���0C|@C��\CYC]Ca3?E?���0�@�
f$�0�d�P�B|@�1 �����!�5(z�O�f+OO;OaO���( �� -�P"�!A!�1�E�S � ���1~Qzр?�ff���O�OfOC �	_[MA8��1_?Z>�!�� DJ(�mUPvX�Isll^�#?���x����<
6b<�߈;܍�<��ê<���<�#^¤�_�AA�+���#$��?ff�f?�?&`�@��.0b�J<?w�\�<bN\�AI �2a
M@to�o gX�O�o�o�o�o �o4XjU�� w���_o�o�o��B��xG@ G@�0�G�� G} t�1���}�����ڏŏ\���BLy3B"�A��T�?��/��I� ?�#	�ϟ-���A��p,�>�P��F�b�I7>�OA @|�����ů��¯���s�A�0��?y5C�M��<>\�?��{���ػ���ѹ�Wy3��fοC 	�CH˿� ��������8�@I���(hA�� �ALffA]���?�$�?��yQӺ°u�����)�	ff��C�#�
��~�g\)Pb�33�C�
������<�p�G��B���L��B�s�����	�RӺH�ۚ�G��!G��W�IYE����C�+�нI���I�5�Hg�MG�3E���RC�j=�
��pI���G���fIV=�E<YDf�Կu�`ߙ� �ߖ��ߺ������� ;�&�K�q�\���� �����������7�"� [�F��j��������� ������!E0i Tf������ �A,eP� t�����/� +//O/:/s/^/�/�/ �/�/�/�/�/? ?9? $?6?o?Z?�?~?�?�?t�?�>(p����o�R��E�5���OOa�3�8�x8OJOa�4MgudO<vOa��VwQ�O�O�4p�+4�] �M�I�O�O __D_2\J��P�RPv^������_�?�_�_�_�_�[R�_o?o*oOouo`o  �@�xo�o�o�o �o�o�_��>,bP{hr���������,���P�>�t���  2 �Fs_�GT�.���Ma�B���,!��C�.�@%�ꏀ��� �2�D�U�����������ǟa�?_���@@Κl��a�a�o�a�p�
 Ο1�C�U� g�y���������ӯ����	��r�� ���`K�D��$P�ARAM_MEN�U ?�E��  �MNUTOOLN�UM[1]]��v�FX�]��A�WEPCR��.$�INCH_RAT�E��SHELL�_CFG.$JO�B_BAS�� �WVWPR.$�CENTER_R�Iϲ��ִAZIM�UTH OPTB���ִELEVATION TC���ִDW��TYP�E SN��ARCLINK_ATڰ?STATUS��7ɿ__VALU��LEP�.$WP_}���gU��|ώ� ��������������0�Y�T�SSREL?_ID  �E�Q��h�USE_PR_OG %c�%U�<��i�CCRTxԐQ�k���_HOST !c�!�����AT�P��+����-��g���_TIMEO�U��g�	�T�GDE�BUGx�c�i�GI�NP_FLMSKĐ��T`����PG�>�  ��n���C�H���+�a�l� T�N߄����������� ��=8J\� ������� "4]Xj|� ������/5/���WORD ?	�c�
 	RS�e	PNH��2gMAI1�p#SU ��|#TEN��3STsYL�s COL
e�1(�/1�TRACE�CTL 1��E�m� tPA |r��&DT Q��E�0� D � �fS��rj+6�5<;�QS0 �Y2�Y2"�Y2��Y0U5U45]45e45m4�5u6��Y2�5W4TW1+6<U4<]4<e4U<m4<u47U47]4�7e47m47�6�3<TF�3<�<9U49]4U9e49m49u44U4U4]44e44m44eFR�39�F�39�<:U4U:]4:e4:m4:u4U6U46]46e46m4I6�F�3:V�3:�; +_=_O_a_s_�_�_�_ �_�_�_�_oo'o9o Ko]ooo�o�o�o�o�o �o�o�o#5GY k}������ ���1�C�U�g�y� ��������ӏ���	�`�-�?�Q��&LE1��z����#  �~�&_UP �;��� ��ñ ��� �� ��$;�ޟ�|�0�  ��)�_DEFSPD ��c�2��  ��T�IN��TROL ���;�8���B�PE_CONFuI����'�Ը�!�0�*LID������	��GRP 1}��) lV��@�j��hs��!A�
D��� D@� Cŀ� @��^� d`���)����0���p"�����C� ´|�^�G�B�����p���𼿦���!>��>�,���7�I�3�� =49X=H�9Nχ�JτϽϨ��� ��f���)���9�_�Jߏ  Dz�Ӎ�� 
 tߵ�d���������� 3��W�B�{�f�x���������)��
V7.10be�ta1Ӗ Aw���6��!���3�?!G�>�\=y�#2�{3�3A!��@����2��8wA���@� A��@�#�B� �����X�����#Ap�"�����dd��$�?����@, �� A|y��33@��#�� Ҿ��7�xߋ� ��ǡ�KNOW_M  �
���SV ]��*�%�� ��������#��"!���Mʣ��-���	ٕ (���ڔ@7X�#�{�3�@{������J ��MRʣ��-�$��`����@/R+��STʡ�1 1�98 4�
Carga_7Too}?�'/���#Pieza ����/�'��ø��/ �/
??.?@?R?d?�? �?�?�?�?�?O�?O@KO*O<O�OW�p'2{,�e4cO  �<�O�Ow 3�O�O�O�O�p'4�O__+_p'5 H_Z_l_~_p'6�_�_�_�_p'7�_ oo$o�p'8AoSoeowop'M�ADw� ��p$O�VLD  ����*}p$PARNUM  ~+s��/�T_SCH�i ���
}wFq�yē�uU�PDFuY���E_CMP_Ow�Ҡ9��'���tER_CHK���ڒ!�
���RS ]��_M�O�`o���_k��E__RES_Gz ���
��J���� ��D� 7�I�h�m�������@�ٟ�o���@Ɍُ ����@(�G�L���GP g��������P��ůʯ ���P��	���@`$� C�H����`c��������V 1�ʅ��e�@]s8��THR�_INR ' dz��d��MASSϛ Z�MN�5�M�ON_QUEUE� �ʅf2�� U��N�UH�NE�nȅ�END�������EXE�Ϥ��pBE����υ�OPTIO��Ǳ���PROGR�AM %h�%�����l��TASK�_I�d��OCFG� �h�\ߏ�D�ATAR����'2p���"�4�F� ��j�|����]�����������INFOR���w�y���e�w� �������������� +=Oas������(�4���� ����ѥpK_��Ѵ��T�G��2�� X,		�R�=���d�'�@�u@}$� `�||�
_EDIT �������WERFL���m#�RGADJ �^�A�  +%?�!�8$
�&���ʅO��,��<|n@T�%�o�/(�M#f�2�Y'�	H��l��f!?#��8A���t$6�*0/2 **�:&2n@?+3G=ʅ�`2[5��1e9΁ �/nB�?S=�=c?u?�? �?�?%O�?�?OOO �O;OMO{OqO�O�O�O �O�O�O�Oi__%_S_ I_[_�__�_�_�_�_ Ao�_�_+o!o3o�oWo io�o�o�o�o�o �o�/Aoew ������]�� �G�=�O�ɏs����� ����5�ߏ���'� ��K�]���������� ɟ�����y�#�5�c� Y�k�寏���ϯůׯ�	��p�l ^����� 9��3��濁�
���I'PREF ��Y*l l 
%IOORITY���!MPDSP�*T��w�UTz��#&OD�UCTw�����&OG� _TG��|����TOEN�T 1�� (�!AF_INE���3�j'!tc�p>�f�!ud�Uߎ�!icmX}ߥ.��XYR#��;�l!)� 31���l ���-��� Y�@�}�d�v����� �������1��U�g�	*��R#�Y)*�/�����l#>��F"1�B37/=<��l$��(��.A{",  �O�Wi{�%���8��@�R�	"!PORT_NUM���l �!_C?ARTREP���;SKSTA�� �LGS0�����{#l Un?othing�s���&�7TEMPG ��ɣ.�[�_a_seiban�/�/</'/`/ K/�/o/�/�/�/�/�/ ?�/&??J?5?n?Y? ~?�?�?�?�?�?�?O �?4OO1OjOUO�OyO �O�O�O�O�O_�O0_ _T_?_x_c_�_�_�_��_�_�_�VERS�I����'` disable����SAVE ����	2670H�771���_�o!`���o�o�߻o 	�hH��0�{��e% N`r�$�=|�o����Gb_�� 1�
��p`�J����� ���1�URGE_�ENB������W�FL�DO�Ƥ�W�,�m���
WRUP�_DELAY ��`�R_HOT %U������~��R_NORMAL�̈��܏1� �SEM�I�6�u�/�QSKKIP�sƺ�sx�_ ���_ޟ��ŝ�3� !�W�i�{�A������� կ�������A�S� e�+�u�������ѿ� ������=�O�a�'� ��sϩϻ��ϓ�������'�9�K�υ�$R�BTIFn�
RC_VTMOU�ջ�i�DCR�sȾ�� �ёB�7șC��MC��g>��k>)P�8���ŝ��<���թ������3y��e�ş�� <
�6b<߈;����>u.�>*?��<���'�� �z��S������ ����	��-�?�Q�c��u��RDIO_T?YPE  �}k����EFPOS1 +1�Oi� x�o
 �h�!E�oi �(��^�� �/A��(�t �H�l���+/ �O/�s//�/�/D/ V/�/�/�/?�/9?�/ ]?�/Z?�?.?�?R?�? v?�?O�?�?�?YODO�}O��OS2 1�����4OnO�OjO_<�O��3 1˨O�O��O_�_o_�_&_S4 1�=_O_a_�_o�o=o�_S5 1� �_�_�_0o�o�o�oPoS6 1�goyo�o��oC.g�oS7 1��o Z��|�zS8 1Б����m�X����SMASK 1ў�� ��Џچ��XNOě�͆����MO�TEp�����4�_CFG �;�������PL_RANG�7�s�u�OWER ��������SM�_DRYPRG �%��%8�����T?ART Ԡ��UME_PRO���ϟJ���_EXEC_ENB  `�{�GSPD#�e�m����|�TDB����R�M����IA_OPOTION�ּ�}�./�MT_��T��9�2��T���c�C�����[�m�����\�i�OBOT__ISOLC��j��g���NAME ���9���OB�_ORD_NUM� ?�����H771  ��B�@B���Bʆ��B��PC_TIM�E��w�xi�S23�2T�1ׯ�̱L�TEACH PENDAN��P���X�7�"@Ma�intenanc�e Cons����ϔ�"��DNo UseX����C��U�g�yߋߏ��NPQO���������oCH_L&��/�悀	���!U�D1:3���R��VgAIL#���ž/�SR  �����o���R_INoTVAL�������ꮅ�V_DAT�A_GRP 2�X����2�D��P�� 1��U�@���x���p� ��������������  H6lZ�~� �����2  VDfhz��� ���/
/,/R/@/ v/d/�/�/�/�/�/�/ �/??<?*?`?N?�? r?�?�?�?�?�?O�? &OO6O8OJO�OnO�O �O�O�O�O�O�O"__�F_/��$SAF_DO_PULS���0���2�pQ`PCANd�����SC�����(�}�����K����R������ J��_
oo.o @oRo�_vo�o�o�o�o��o����kb2$�dڍd�dqF�s�� @n�@Rd�v~(y� ��t_�_ @�T���������T D���-�?�Q�c� u���������Ϗ�� ��)�;�M��߱�:u/�������o����;�o�����p���
�?t��Dia�la��Q��  � � Ϻ�QlaR��Q;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟπ����������ߕ�� ;4�F�X�j�|ߎߠ� ������e����&� 8�J�\�n������r0���(����� ��+�=�O�a�s��� ������������ '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�ߝ/�/�/�/�/ �/	??-?������kb m??�?�?�?�?�?�? �?O!O3OAITOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o:o��c��Eo�o�o �o�o�o�o�o $ 6HZl~��Jj�oo�������-��_�	12�345678��h!B!ܺ[4��m`��V�h� z�������ԏ�� no�!�3�E�W�i�{� ������ß՟���� �/�@���c�u����� ����ϯ����)� ;�M�_�q���B�T��� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/���S�e�w�� ������������ +�=�O�a�s���D�� ��������'9 K]o����� ����#5GY k}������ �//1/�U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?NcG��?�?K/�?�?�O �Cz  B}pKj   �]hu2abG�} Lh�
]G�  	�Nb2�?�O�O�O�O�KK>�9DFo�<�wO _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro_�o�o�o �o�o�o&8J \n��������I.B�1kACB�<-��$SCR�_GRP 1���8� � �� �.A �>E	 b��j�{�t� �1���,G������܏�M�M@قD��W�N���ً�L�	M-10iA/�7L 12345_67890m@P�; 8m@MTW�_�&.C
Z����\�]KSB��_j�.FY���Y��Cف�Ax�����	SJ�"�4�F�X�.D?��H�j��n�Y�������ǯٯ���o.A�����A���3�p���B�'@Ɛ��������A8@�� C @.@ʵ���?�@�򵆲H'@�ݺ��F?@ F�`-�5� ,�Y�D�}�hύϳϞ� ������~�ʱ��&��#�5�G�B�U��ϛ� �߿ߪ��������� =�(�a�L���O���ŏ����>G_@��
�x.B�ʱ=m��DȰ��@ʰJ�'@�`�Z������?��.DCA����������A��.A �������BN`/ (� �����}����.F9�EL�_DEFAULT�  Ô���.@HOT�STR&��8�EM�IPOWERFL�  E2`W�FDO' tR�VENT 1����s�Q L!�DUM_EIP�,H�j!AF�_INE&�.D!'FT�.�>/9!��c/ �-/�/�!RPC_MAIN�/m(�y/�/�#'VIS�/l)��/"?o!TP0PU?��d?n?!
PM�ON_PROXYo?�e]?�?52�?��f�?O!RDMO_SRVO�g�?�RO!R��nO�h,AO�O!
� M�?��i�O�O!RLSgYNC�O��8�O>6_!ROS�]\��4%_�_!
CE>70MTCOM�_��kq_�_!	�RCO�NS�_�l�_o!}�RWASRC!O��m	ofo!�RUSBgo�nUo�oQ/ �oC�o�o�o$�oH�l3�RVI�CE_KL ?%�� (%SVCPRG1����u2���p3���p4/�4��p5W�\��p6����p7�����pH{���|9�����t iO$��q�L��q�t� �q!����qI�ğ�qq� ��q����q��<��q �d��q����q:��� �qb�ܯ�q����q�� ,��qڟT��q�|��q *����qR�̿�qz��� �q����ʯ��r�p ��pgϬ��q���Ͽ� ������@�+�d�v� aߚ߅߾ߩ������ ���<�'�`�K��o� ������������&� �J�5�n�Y������� ����������4F 1jU�y�������0�z_D�EV ���MC:o�4���JGRP 2��o��pbx 	� 
 ,�8�o�� / ��6//Z/A/~/�/ w/�/�/�/�/�/?�/ 2?D?�h??�?�?�? �?�?�?�?�?OO@O 'O9OvO]O�O�O�O�O �O�OK?�O*_�ON_5_ r_�_k_�_�_�_�_�_ o�_&o8oo\oCo�o goyo�o_�o�o�o �o4-jQ�u �������� B�)�f�x��o��S��� ҏ����ݏ�,��P� 7�t�[�m�����Ο�� ���(���^�� ��i�������ܯï � ���6��Z�l�S��� w��������A�� � �D�+�h�O�aϞυ� �ϩ���������@� R�9�v�]ߚ߬���� �������*��N�`� G��k�������� ���&�8��\���Q� ��I����������� ��4F-jQ�� ������id �i	U@�yd���)%�x��q����! �%/,'/L/:/p/ ^/�/�)��/
)�/�/ �/??(?*?<?r?�/ �?�/b?�?�?�?�?O O$Oz?�?qO�?JO�O �O�O�O�O�O_RO7_ vO _j_�Oz_�_�_�_ �_�_*_oN_�_Bo0o foTovo�o�o�oo�o &o�o>,bP r��o��o��� ��:�(�^������ N�p�J����܏� � 6�x�]���&���~��� �����؟�P�5�t� ��h�V���z������� �(��L�֯@�.�d� R���v������$� ����<�*�`�Nτ� ƿ���t���p���� �8�&�\ߞσ���L� �ߤ����������4� v�[��$��|��� �������N�3�r��� f�T���x�������� ��������,bP �t����� �(^L�� ��r�� /�/ /$/Z/��/�J/�/ �/�/�/�/�/?b/�/ Y?�/2?�?z?�?�?�? �?�?:?O^?�?RO�? bO�OvO�O�O�OO�O 6O�O*__N_<_^_�_ r_�_�O�__�_o�_ &ooJo8oZo�o�_�o �_po�o�o�o�o" F�om6X2� �����`E�� �x�f�������ҏ�� ��8��\��P�>�t� b�������Ο���4� ��(��L�:�p�^��� ֟��ͯ��� ��$� �H�6�l�����ү\� ƿX�ֿ��� ��D� ��kϪ�4Ϟό��ϰ� �������^�C߂�� v�dߚ߈߾߬����� 6��Z���N�<�r�`� ������������� ���J�8�n�\����� ������������� F4j�����Z� �����B� i�2����� ��JpA/�/t/ b/�/�/�/�/�/"/? F/�/:?�/J?p?^?�? �?�?�/�??�?O O 6O$OFOlOZO�O�?�O �?�O�O�O_�O2_ _ B_h_�O�_�OX_�_�_ �_�_
o�_.op_Uogo o@oo�o�o�o�o�o Ho-lo�o`Np r���� �D �8�&�\�J�l�n��� ���ݏ������4� "�X�F�h���䏵�� ���֟���0��T� ��{���D���@���� ү���,�n�S���� ��t��������ο� F�+�j���^�Lς�p� �ϔ϶�����B��� 6�$�Z�H�~�lߢ��� ���ߒߴߎ���2� � V�D�z�ߡ���j��� ��������.��R��� y���B����������� ����*l�Q��� r�����2X )h\J�n� ��
�.�"/� 2/X/F/|/j/�/��/ /�/�/�/??.?T? B?x?�/�?�/h?�?�? �?�?OO*OPO�?wO �?@O�O�O�O�O�O�O _XO=_O__(__p_ �_�_�_�_�_0_oT_ �_Ho6oXoZolo�o�o �oo�o,o�o D 2TVh��o� ����
�@�.�P� �����v�Џ��� ���<�~�c���,� ��(���̟���ޟ� V�;�z��n�\����� ��ȯ���.��R�ܯ F�4�j�X���|���Ŀ ��*�����B�0� f�Tϊ�̿����zϜ� v�����>�,�bߤ� ����R߼ߪ������� ��:�|�a��*�� �����������T� 9�x��l�Z���~��� �����@�P���D 2hV�z���� �
�@.d R����x�� /�/</*/`/��/ �P/�/�/�/�/?�/ ?8?z/_?�/(?�?�? �?�?�?�?�?@?%O7O �?O�?XO�O|O�O�O �OO�O<O�O0__@_ B_T_�_x_�_�O�__ �_o�_,oo<o>oPo �o�_�o�_vo�o�o �o(8�o�o��o ^���� ��$� fK���~������ ��؏Ə��>�#�b�� V�D�z�h�������ԟ ���:�ğ.��R�@� v�d������ӯ��� ���*��N�<�r��� ����b���^�̿�� &��Jό�qϰ�:Ϥ� �ϴ϶�������"�d� I߈��|�jߠߎ߰� ������<�!�`���T� B�x�f�����(� ��8���,��P�>�t� b������������� (L:p��� ��`�����$ H�o�8�� ����� /bG/ �/z/h/�/�/�/�/ �/(/??�/�/�/@? v?d?�?�?�? ?�?$?�'1�$SERV_MAIL  .5�$@�
HOUTP�UTH�
HRV 2�6  '@ (�1�?�O�DTOP10 2}�ZI d *? �O�O�O�O	__-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m�����5�EYPE�:L(EFZN_CF�G �5�'C'4IB�xGRP �2��w�q ,B�   A?�'1D;� B@��  �B4'3RB2�1�FHELL�r!�5�vm@nO���>�;%RSR���� ʏ��'��K�6�o� Z�l�����ɟ���؟��#�5��  ���5�c�u�C��� '0}�����'8K��2'0d�����j�H�K 1�x�  ���$��H�q�l�~� ������ƿؿ����� �I�D�V�h�d�OM�M �x���i�FTOV_ENBD�bA�u��OW_RE�G_UI��BIM�IOFWDL���x��B��WAIT��A٩IE8�4@��aD�2�TIM�����l�VA@C��_U�NIT�ã��yLC���TRY���u�@MON_ALI_AS ?e��i@he�?'�9�K�]�%: ������o����� ��0���T�f�x��� ��G����������� ,>Pbs�� ��y�(: �^p���Q� �� //�6/H/Z/ l//�/�/�/�/�/�/ �/? ?2?D?�/h?z? �?�?�?[?�?�?�?
O �?O@OROdOvO!O�O �O�O�O�O�O__*_ <_N_�Or_�_�_�_�_ e_�_�_oo�_8oJo \ono�o+o�o�o�o�o �o�o"4FX |���]��� ���B�T�f�x��� 5�����ҏ������ ,�>�P�b�������� ��g������(�ӟ L�^�p�����?���ʯ ܯ� ���$�6�H�Z� �k�������ƿq�� ��� �2�ݿV�h�z� �Ϟ�I���������
� ��.�@�R�d�߈ߚ� �߾���{�����*��<����$SMON�_DEFPROG &���f�� &*SYSTEM*C����R S�RECALL ?}f�� ( �}3x�copy fr:�\*.* vir�t:\tmpba�ck��=>192�.168.56.�1:14432 `��������}4��a��������������}8��s:ord�erfil.da�tP�b�x�	-}=/��mdb:M��� �������:���T� f�w,?��� u��������Xs //(/;M�q�/ �/�/�L^� ?? $?7I�/m~?�?�? ��P/��?O O3/ E/�?i/zO�O�O�/�/ V?�/yO
__�OA?�O �O�O�_�_�_�?�?ZO uOoo*o=O�_aO�_ �o�o�o�ON_`_�O &9_�o�oo_�� ��_�_Ro�_��"� 5oGo�ko|������o �oX�o����1C ԏg������/��� \�w���,�?�ڟc� ����������P�]�� ��(�;�̯ޯq��� ������˟T�� �� $�7�I��m�~ϐϢ� ��ǯZ����� �3� E���i�zߌߞ߱�ÿ տc�y�
���A��� e��߈����R�_� ����*�=�����s� ����������V��� &9�M���o�� �����\����" 5�G��k�|���� ��Ne�//1C��g��/�/�.�$�SNPX_ASG 2�����!��  �0�%��/�/  �?��&PARAM� ��%�! W�	�+P����I4�� OF�T_KB_CFG�  ��%�#OP�IN_SIM  �+D2�?�?�?��3� RVNORDY_DO  N5�v5�2QSTP_DSB�>D2"O�+�SR ��) G� &H:eO��&�TOP_ON_E�RR�?�FPTN ��%�@��C�BRING_P�RM�O�2VCNT?_GP 2��%F1� x 	O_�`_@_+_d_�'VD�@�RP 1�9G0 UQ�1G_�_�_�_�_�_ ooo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�`�]�o��������� ɏۏ���&�#�5�G� Y�k�}�������ş� �����1�C�U�g� y���������ӯ��� 	��-�?�Q�x�u��� ������Ͽ���� >�;�M�_�qσϕϧ� ���������%�7� I�[�m�ߑߣ����� �������!�3�E�W� i����������� ����/�V�S�e�w� ���������������+=Oas}RP�RG_COUNT�k6�B�	ENB��O�M�m4�_U�PD 1�HKT  
��-? hcu����� ��//@/;/M/_/ �/�/�/�/�/�/�/�/ ??%?7?`?[?m?? �?�?�?�?�?�?�?O 8O3OEOWO�O{O�O�O �O�O�O�O___/_ X_S_e_w_�_�_�_�_ �_�_�_o0o+o=oOo xoso�o�o�o�o�o�o 'PK]o �������� (�#�5�G�p�k�}���𸏳�ŏ�_INF�O 1�	�  ��� �,��P�;�@����>P`>�����W��A���BU?�N�������´��YS�DEBUG� 
��׀d�	��SP_PwASS�B?̛�LOG �	]  ׀׈��  ��ׁUD1:\�����_MPC��	z����	5��� 	Z�SAV ���B��!�9�ׅ@�SV���TEM_TIM�E 1��� 0  ���Պ9��SKMEOM  	�!�  ׂ%H�����.ׄ� @׀��ׁ4�ׁ"ׅ5��� AJ�p p̼�0�*׃HʰׁB�nϐ�ϒϤ��^���V W��κ˳��
�� .�@�R�d�v߈ߚ߬��������R���%� 7�I�[�m����� ���������!�3�E��W�i��T1SVGgUNS�'���~�ASK_OPTION� 	����_DIې����BC2_GRP 2�	�+���k�˰�C�׉A��*��*׀V9.00�55 C1/31�/2017 Ac w�11M���_ACC_T���X-$tLEN_1  �2��EL_RA��� �$��W_AXISV�F1tI�2��MOVE����E�RTIA  � 	$D�TORgQUEs�DE���LACEMNT��t ��V� MA�XAATCV8HiTRQh�^STAT�L�J_��M��� J_MOD�;$D� ��2�P�!6� JK&VK�1!4�1!3##J0F$5#�JJ=#JJE#AAAL5#k =#k e&4f%5��N1�� [�E�L� _NUM���oCFGw� ` $GRO�UPDSK�B_CONFLIC��� REQUIRE�D����p�$T2 -1q 6o�SG��w \ $ENABL��$APPR#0C�L�
$OPEN�j8CLOSEy:SC_M��� �9
o�PARA�  �b0MCD��^�4_MGN�3C���AV�9�C�7BR�K�9NOLD�6S�HORTMO_L!I�!#GM�5J,@DPm$#=##E##�#�#�##6ZE7ZE8�!�oM4�  2���G��CPATH�G�A�C�AР�C�020� CN�Tj0A^2#Gk2�1I�NsUC� �3PC��UM<XY� 0�CQYP_E� ^Z� �^ZE ^PPAYLO�AGJ2L_UP�R_AN1�SLW�[�Q�Y�Q�5R_F�2LSHR��TL�O�T2Q�W@S�W@SACRL_�0U#`,WܑT�HVAm3$yH�2QbFLEXm3��o J��w MPW2B_� �!� M_FTM��d�?RESERVjQ�g̡jE!mas :���g�d������F1 �aHu\w���+�rE5GYk} ����c����� $pp����
/�a*	T��a�X<pi�%�t �x(%1�
�4/F/X/j  n%w%e%�%�/�/�/�)��lb�$ � ��/�/?�UPDA1Tuv1�EL�p+��F�&8J20-0JE�
@CTR,QpqTN�pFC�7HAND�_VB�rmaOPnL5 $ՀF2�6��3]�COMP_S�W�aC3�6	� '$$M�P�9R�3���	A��p��B"�A_��R�6D<��=A�<A��<AKAKJ��;D��<DKDKP�@GR�7�ST�7�	I�NHDY�Ph0�6 +�R��Pu �W�a�W�Q@�W'��"p�EPbE kEtE}E�E�E�E�B�2JL5
 ��d�B� �q�Ŝ1��AS�YMUh`��V	p#�"]�Q'__SH�" 1WKT5M7Ի�U_g_y_�_�SJ�\U@�Z����\�Y�t_VI���|�3$�V_UNI�S8�Z��QJ %Q��Q� �\U�eb��m�'i U@6oHo���^dfc� ��TO0HR_T\2�����a1DI@ƃO&����@��#��
Y�I<�A�1@SS�vp�a�a��pS��`�p	� � � ̡M�E�q��|���c�T�PT��ؐ�@��� ��$Y0�Щ����T����! $DU�MMY1b�$P�S_spRF5p! u$���0FLA� �YPŃ��$GLB_T��4���`1l`�pt�B� XXW07M1ST�q-0�SBRPM21_�Vg�T$SV_E�R�PO��z�CL�N zA�pOV��G�L�EW�! 4\� ��$Y/rZ/r!W� �QȣA}�<Rt���U� ՀyN� ��$GI���}$� q�� �! L� \��}$F��E �NEAR�pNzsF�g�pTANCzr�?��JOG)pK@�   $JOINT��p��MSET�!  "EM�q�S��0�4��!� �qpU�q?�-0LOCK_FO�Pӡ"�oBGLVw�GL(TEST_XMm0N�EMP�g�5"L�$U�`��2,1�[!&"Ϡ [!|CE� )| _ $KAR'�M(�TPDRA� �$��VEC�`�&�IU�[!{CHE TO�OL<s�#V;tREN� IS3�e�"6��NppACH�h��!1OP����29��� �I]2  @$R�AIL_BOXEz�� ROBO,$�?��HOWWA�RYaK1��1ROLMq5ב4�2�90�@p�@O_F�!C �A� 	1�A�W �R� O�b�2�4p��07�OU�bW%��M�'���$PIP-&N À�"92	1�p[!�0�`?CORDED h���0y�P�Oc� � D 3 OB �Q� nG]A��2 ]B܍�S�SYS]AADqRR���TCH��  ,ՀENT�aA!_�D����a WAVWVA~� � � ���PREV_R�Tt�$EDIT�VVSHWR�Pf.P�r��D����aETq$HECAD����_P��S�KE���CPSP]DvVJMPz@L�2ڠR�p>�e@~a��FI6 SR�C��N�E� S���TICK�<sF�M��A�SH=N\ @g@�Q�~Q_GPf06�`gSTY�B1LON� �T	b�� tk 

PG�E%$�A�=f SH�!$@G����P�P)�fSQU� /u �TERC��/q��S� r � À����!5�O���F2pIZ!��PRO@+r�Q�0P9U�;u_DOl�@�XS�K�AXI4Zp�3`!UR ��s@S�R0�P�Fá!�_� �BET�rP
"v@�%Y`F�Z`A��C��*3$3j��{SR��l�` �$�����(�"�� -��;��K�\�m�\� }�\���n�����n��� �������C����p�ߪ߼��SSC6 �   h� DS�`�!��SPM���A	T{�#�<q�P�R��ADDRES�#B�PSHIF�R _W2CHR��AIU �ڑ�TUU I� �!�2CUSTOT�t�1V�IA�"�BP(��s��
5*
7�qV�1Kq^ # \�P�H�Y`*��a�g�C����b�r9�F�g��TXSCREE_B�$�uaTINA�&���A�q����% T�Q� r�A �q �hq�Bhr�PRROV���@pP ��t�QUE�T& �����A S��ARSyM�P^wUNEX�`�q��S_���@� ������@ӜqC�m��� 2%��UE���'G�Զ+pGM�T��Ls�wq� O���`BBL_0W���^ ( �Y`1�O�=�LE̒H�Q0� �G�RIGHQ�B�RD�CKGR��y�TEX�pz�u�WIDTH3;Pr�,1�!�UI�0EY��]) d�� P�=b90'qB�ACK;a�ū��FOFA��LAB�F�?(��I0�$URW1,л ����}H'� * 8��B�_^QڒOҎ�R� @�$37���<�OӑJ^ +`�r�U]�r��R
"|1LUM�Ӝv��ERVA9�P�k��,���pGE�0�R�p�)gPLP$���rE�`M�)�lQ��m��0�5�6
�7�8���b��&pPk{���1�S��+��USR�'- <�P��U��FO��PRI��qm#0����TRI}P51m�UN.�
?�.~`.�Uc1�_u�S!�p�` /�Jҹ�*qG f`T0�0;�ۑE�OS��Z�AR�p-�1��!]0�@����d�0R"U��]1��������e1�OFF+ ^ 2b z��O  10� ���"1� GU�AP�!�=8�G��SU1Bb� 0�RT���ta3b��0
sOR0N�RAU��T�	��G�VC>�84G� /2^A�cb$���a3�C�0�D�RIVv�q_V�`2P�D��MY_UBY���`f�� �e9��`ҠLQo�!~P_Sz@jt A{�BMD�$�PDEY�CEX�E�&�`_MU�PXD����US{�� ��� Ѡ�b����9��aG̀PAgCIN�Q�`RGMp %#"��#"��#"���CREd�Б�!�2��#"�05 �0TARG)P��h �@�	Rq�06����iq���m	�XqRE�SMW _A!�p�)pO��AԐ�#�EE��UL`1�p��V�HKQb7`�*`�`�� �%3EA�P�/7WORQ��%�%MwRCV�8 ���UO]`MQ�C��	l28��e#l2REFǎ6 u6`1� ���s� ��q:��1�:�1�;�5u6?_CRC0;HI;��S����5�a�A��l"�9 �.b�����`��:�`OUg`"f�O 4~%<�2R�a$��}�*p�P6��t<��RK{pSUL���7��COe�f�8��@JS
�SXQV ~�V��S�@Lz9U`�9U~�EW����>�T:| +���qzՠ ��CACH5cLO�1�T�Q��Yq����cC_LIMI͓FR�XTt��VVK�$HOQ�mb�PC'OMM�m�O[�g`H��уDd�VPb"$�@Kb_vUdZ Phl�PPhWA�UMPujWFAI�PG!4�P�AD�i�IMRE�D�bZgGPs�����ASYNBUF�VRTD�etZa6��OLՐD_��uuW��P�ETU��PQ� �eECCUU(VEM? �Ugr�WVIRC�au�cl�>q_DELAZ#�X8��kAGyR�GXYZ�����W�!�s���pT� �.��r�;����LAS��H�1pQc�G�a{�<�ҾQS�`�VN<�,�_VLEXEwU=��d�����^cFLv�I��cFI!p��@~��"3p�r��t">��d�\D���b.H�ORD������T�B5�?Š��T���XO���Ґ S9F��U�@  Ǡ��Q�URR3<�MF�A���J��f���a�B�$�N�LIN��m��MW�0XSK1��CJ��%�F@K��H��HOuLс�!XVR
��D�	�T_OVR~т
�ZABCzAEz"�׃��V1ZD �
�F�DBGLV�OcL5���ZMPCFzGJ�k�(��}�DLN䐜0
qj��{H ���xa/0��CMCM }COcCART_����$P_�� $JݣפD@a���`�s���sМ2UX�q��UXE�'��q����J�0�B�0�R�<�A�I }�\��U0~�Y��D4� �JJ�R�`���pH!Ek���%� ��������mDK � �1��18�s�EAK|�7@K_SHIP�,Vp��RVypFv�2#��C?�آ͡�D2���>���BIf�5eD�v�TRACEa�V|�q}�SPHER��L ,�@��п⹿�$TBCs� ������?�  `�ɗ �����`���	�O�:� L߅�pߩߔ��߸��� ���'��K�6�o�Z� ��~��������� ��5� �Y�D�}�����{���|�����j��� %I4m���ő��a����� �'79K� o������� #//G/5/k/Y/�/}/ �/�/�/�/�(���/? -???Q?�/u?c?�?�? �?�?�?�?�?OO;O )O_OMOoOqO�O�O�O �O�O_�O%__5_[_ I__m_�_�_�_�_�_ �_�_!ooEo�/]ooo �o�o�o/o�o�o�o �o/AS!we� �������� =�+�a�O���s����� ��ߏ͏��'��7� 9�K���o���[o��ϟ ������5�#�E�k� Y���������ׯů�� ���/�1�C�y�g� ���������ӿ��� 	�?�-�c�Qχ�uϗ� �ϫ�����߻��/� M�_�q��ϕ߃ߥ��� ��������7�%�[� I��m�������� ����!��E�3�U�{� i��������������� ��A/e�}� ���O��+ OasA��� �����/9/'/ ]/K/�/o/�/�/�/�/ �/�/�/#??G?5?W? Y?k?�?�?�?{�?�? OO1O�?UOCOeO�O yO�O�O�O�O�O�O_ 	_?_-_O_Q_c_�_�_ �_�_�_�_o�_o;o )o_oMo�oqo�o�o�o �o�o�o%�?=O m���������v-��$TB�CSG_GRP �2�u��  �-� 
 ?�  X�j�T� ��x��������ҏ���1�8��G�d�, �M�?-�	 �HCA�����i��CS�B�P�����]�>���ͱ�u�Г�۝B���333���Bl"{����#�Aʐ��fffA��5�C��#�%��s�?�� ��N�~�Y���A-��ӧš����@ƯP�� 4����_�|�G�Y����Ŀӻ�����	V�3.00P�	mt7���*��,���ݶY��@f�f-� -�H�� �U�'�V�  �����'ϖϟ�1�J2�8�?��ϫ�CFoG �uI�Y L������k�*��*�P�^�� ^߄�oߨߓ��߷��� ������J�5�n�Y� ��}���������� ��4��X�C�|�g�y� ����������P�jp );��nY~� �����"4 FjU�y�� -������/C/ 1/g/U/�/y/�/�/�/ �/�/	?�/-??Q??? a?c?u?�?�?�?�?�? �?OO'OMO;OqO_O �O�Og�O�O{O�O_ _7_%_[_I__m_�_ �_�_�_�_�_�_�_3o !oWoio{o�oGo�o�o �o�o�o�o�o/S Awe����� ����=�+�M�O� a���������ߏ͏� ��9��OQ�c�u�� ��������ɟ���#� �G�Y�k�}�;����� ů��կ����ٯ/� U�C�y�g��������� ѿӿ��	�?�-�c� Qχ�uϗϽϫ����� ���)��9�;�M߃� qߧߕ����߇���� ����I�7�m�[��� ������������ E�3�i�W��������� }�������A/ eS�w���� ��+O=s a������� //%/'/9/o/�߇/ �/�/U/�/�/�/?�/ 5?#?Y?G?}?�?�?�? q?�?�?�?�?O1OCO UOO!O�OyO�O�O�O �O�O�O_-__Q_?_ u_c_�_�_�_�_�_�_ �_oo;o)o_oMooo �o�o�o�o�o�o �/+=�/�om� ������!�3� E���{�i�����Ï Տ�������-�/� A�w�e���������� џ���=�+�a�O� ��s�������߯ͯ� �'��K�9�[���o� ��QϿΉ����� �G�5�k�YϏ�}ϳ� �����ϧ������ 1�g�yߋߝ�W��߯� ����	�����-�c� Q��u�������� ���)��M�;�q�_� �������������� 7I�as�/ �������3 !Wi{�K��p����   �## #&7/#"��$TBJOP_G�RP 2���  ?��#&	O"V#
],����� ��� =r%  Ȯ� � �� �#$� @ n"	 ��CA��&��S�C��_#%n!�"G;��"k��/;�=�CS�??��?�-0,0?CR  B4�'F?xQ7�/�/?333�2�Y-0�?�:;��v�'2�1�041*90��=?�?90��7C� � D�!�,� BL���O%K:�Z��Bl  @pI@�^� s33C�1 �?�nO  AЁG�2�qG�&0A0E�O�J;����A?�ff@,\@�1C�a0zqO�O��@���U�O�$f�ff7R0_B^;xCsQ?ٽ40@�O�_�{F�X_Q\LU�_�V:'�t-�Q/B�1@�O o!h�&4h+oaGSo=o Koyo�o�o?o�o�o�o �o	:�oYs]Pk��]4�#&`�q��%	V3.00�t#mt7H@�*��s$!#�.� �E��qE����E�]\E�H�FP=F�{�F*HfF@D��FW�3Fp?�F�MF����F�MF���F�şF���F�=F����G�G.�?�CW�RD3l�)D��E"���Ex�
E���E�,)Fd�RFBFHFn�� F��F���MF�ɽF�,�
GlGg�!G)�G=���GS5�Gi���;��
;�Uo�|& : @_zQ-/�%�#&)��?�0�&[�B-ESTPARS  (�h L#HR~�ABL�E 1]) $G�##i�>� � �
i�i�i�"'*!i�	i�
i�i���#!Ui�i�i���'RDI��g!��ɟ ۟����y�O����@������ӯ宙�S�e# C�����ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ���������B- ~���f"��=�&�8�J� \���,�>�P�b���~#�NUM  ��g!� +  ���t���_CFG ����!@O IMEBF_TT��0��e#��N�VE80t��O�d�N�R 1��� 8 �#"d �� �H�  �� ����������'�9� K�]�o����������� ����6#lGYo}��ANӹ��V;MD��� 8%7IV_I]o�IINT��IT��� Bf�	//��
_TC=/O/I$0��w/�/�RQ�/�/R��_�{�@��{�MI_CHANZ�� �� (3DBGL�VLZ���z�+0E�THERAD ?U��~0�)��/��/�?�?s�+0ROUmTx�!
�!�4��?�<SNMASK�s8��1255.�9E�7OIO[O�{�O�OLOFS_DI��%]9ORQC?TRL ���*��MT�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo-l�OPo�?otox�PE_DE�TAIQ8�JPGL�_CONFIG ��ᄀ/�cell/$CID$/grp1xo@�o $6죀�? as����J� ���'�9��]�o� ��������F�X���� �#�5�G�֏k�}��� ����şT������ 1�C�ҟ�y���������ӯG�}h�	��-��?�Q�c���eo��j�� g���ҿ�����a� >�P�b�tφϘ�'ϼ� ��������(߷�L� ^�p߂ߔߦ�5����� �� ��$��H�Z�l� ~����C������� � �2���V�h�z��� ����?�������
 .@��dv��� �M��*< �`r�������`�User� View �i}�}1234567890�/!/3/E/`W/_$� �c/���2�\�/�/�/�/	??z/�/�3�/i?{?��?�?�?�?"?�?�.4 X?O/OAOSOeOwO�?�O�.5O�O�O�O_ _+_�OL_�.6�O�_ �_�_�_�_�_>_ o�.7t_9oKo]ooo�o�o�_�o�.8(o�o�o�#5G�ohnr �lCamera��o�������E�1�C�U� �o���������ɏ�I  �v�)��+�=� O�a�s����������ߟ���'�9�`� �vW9П��������ͯ ߯����'�r�K�]� o�������L�^�I<� ���'�9�K��o� �ϓ�޿���������� ߸�^�勪�_�q߃� �ߧ߹�`������L� %�7�I�[�m��&߈u sY����������#� ��G�Y�k�������� ��������^�'i��5 GYk}�6��� �"�1CU ��^��i����� ���/1/C/�g/�y/�/�/�/�/hz9 M/??&?8?J?\?/ m?�?�?K/�?�?�?�?PO"O4O�j	�u0�? oO�O�O�O�O�Op?�O �O_�?5_G_Y_k_}_ �_6OHO�p�{3_�_�_ oo0oBo�Ofoxo�o �_�o�o�o�o�o�_ �u���oTfx�� �Uo���A�,� >�P�b�t�UEh�� ��ҏ������>� P�b�����������Ο ������Իw�,�>�P� b�t���-�����ί� ���(�:�L�󟙅 @�㯘�����ο�� ���(�:υ�^�pς� �Ϧϸ�_�����O�� �(�:�L�^�ςߔ� ���������� ��$���  ��S�e� w�����������<��   )�1� O�a�s����������� ����'9K] o������� �#5GYk} �������/ /1/C/U/g/y/�/��  
��(  }�G�( 	 �/ �/�/�/�/??=?+? M?O?a?�?�?�?�?�?:�*9� �s�$O 6OHO��lO~O�O�O�O �O��O�O__[O8_ J_\_n_�_�_�O�_�_ �_!_�_o"o4oFoXo �_|o�o�o�_�o�o�o �oeowoTfx �o������= �,�>��b�t����� ���������K�(� :�L�^�p���ɏۏ�� ʟܟ#� ��$�6�H� Z���~������Ưد ���� �g�D�V�h� ��������¿Կ�-� ?��.�@χ�d�vψ� �ϬϾ�������M� *�<�N�`�r߄��Ϩ� ���������&�8� J�ߣ߀������� �������"�i�F�X� j�������������� /�0w�Tfx�������0@  ������ ���#frh:\�tpgl\rob�ots\m10i�a;_7l.xml�_q����`���/.��/ 8/J/\/n/�/�/�/�/ �/�/�/�//?4?F? X?j?|?�?�?�?�?�? �?�??O0OBOTOfO xO�O�O�O�O�O�O�O O_,_>_P_b_t_�_ �_�_�_�_�_�_	_o (o:oLo^opo�o�o�o �o�o�o�oo�o$6 HZl~���� ��� �2�D�V� h�z�������ԏ�t��P ��%<< #?���;���3�U��� i����������՟� 	�7��?�m�S�e��������������$T�PGL_OUTP�UT / �#�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϠϲ�����#�����2345678901���� 1�C�U�]����τߖ� �ߺ�����v����&�8�J�\���}f��� ������n����0� B�T�f���t������� ����|���,>P b������� �� (:L^p ~������ �$/6/H/Z/l/~// �/�/�/�/�/�/�/
? 2?D?V?h?z??$?�? �?�?�?�?
O�?O@O ROdOvO�O O�O�O�O �O�O_�O��}�<_@N_`_r_�_�_�]@���_�_#� ( 	 ��o o6o$oZo Ho~olo�o�o�o�o�o �o�o D2Tz h�������@�
�@�.�d��Ƹ� 2�l�������ҏ䏾� ���ʅ�K�]���i� ��m��ɟ۟9�ߟ� ����G�Y�3�}���� w�ů_�������1� C���+�y���%����� ��Ϳ��U�g�-�?�ٿ G�u�O�aϫϽ���� �ύ���)���_�q� ��yߧ�Aߓ������� �%���[�m��� ��}����7����!� ��E�W�1�C������� ����o�������A S��W�#u�� ��e�=�) s�_���� /�'/9//E/o/� ��/�/Q/�/�/�/�/ #?5?�/Y?k??W?�?�{?�?�?�?{��$T�POFF_LIM� ���@|�y��ABN_SV@�  �TJP_�MON x�)D�@�@2�UA�STRTCHK �x�F9_"BVTCOMPAT/H��AFVWVAR �OM�H3D ��O �O@bB�A_DEFPRO�G %~I%�MAIN_MANIPULACIJ@�R_"B_DISP�LAY@~N$RIN�ST_MSK  �v\ `ZINU�SETP�O$RLCK��\[QUICKM�EN�_fTSCRE��Px��BtpscfT�Q`iB�,`_0iST�JIR�ACE_CFG �OI�D@	��D
?�whHNL� 23ZX��a�K  	R�o�o�o);�M_zyeITEM �2�k �%$�12345678�90��u  =<����s  !��{P�?��C� `����������0� ��T��x�$�J�Џ�� ҏ������,�؟�� �t�4�������6��� ����į(�ЯL�^�p� ��B���f�x�ܯ�� � �ۿ6���Z��,ϐ� Bϴ�Ϗ�꿪�Ϻ� ����V���zόϞ�� ��nߔߦ�
���.�@� R����߈�H�Z��f� ���߽����<���� r�$����q������ ����H�8�J�\�v��� ����Pv���� "4�X*<� H���l�� �T�x�S/�n/ ��/�//�/,/~/? b/"?�/2?X?j?�/v? �/??�?:?�?OO �?BO�?�?�?NOfO O �O�O6O�OZOlO5_�O P_�Ot_�_�O�__ _��_udS�b�o�Zψ  jr�Z 8�aEo<Y
 Roxo�_o�ojUD1:�\�l�� aR_G�RP 1�{?� 	 @EP�o {�o&J8n\~�~p��zhq�o��<��u?�  �� �>�,�b�P���t��� ������Ώ��(��0L�:�\���	�U������SSCB 2 
k ������*�<�N�`�r����\U�TORIAL �!
k�oϯ�WV_C�ONFIG "�
m�aBo�o.�ޭOUTPUT #
i���:�~��� ����ƿؿ���� � 2�D�V��k�~ϐϢ� ����������� �2� D�V�g�zߌߞ߰��� ������
��.�@�R� c�v��������� ����*�<�N�`�q� �������������� &8J\m��� ������" 4FXi|��� ����//0/B/ T/f/w�/�/�/�/�/ �/�/??,?>?P?b? s/�?�?�?�?�?�?�? OO(O:OLO^Oo?�O �O�O�O�O�O�O __ $_6_H_Z_l_��i� �_�_�_�_�_oo(o :oLo^opo�ouO�o�o �o�o�o $6H Zl~�o���� ��� �2�D�V�h� z������ԏ��� 
��.�@�R�d�v��� ������П����� *�<�N�`�r������� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϟ��������� ����0�B�T�f�x� �ߛϮ���������� �,�>�P�b�t��� �߼���������(��:�L�^�p�����wX���������� ���_&8J\n ��������� "4FXj|� ������/ 0/B/T/f/x/�/�/�/ �/�/�/�//?,?>? P?b?t?�?�?�?�?�? �?�??O(O:OLO^O pO�O�O�O�O�O�O�O  _O$_6_H_Z_l_~_ �_�_�_�_�_�_�__  o2oDoVohozo�o�o �o�o�o�o�o	o. @Rdv���� ����*�<�N� `�r���������̏ޏ ����&�8�J�\�n� ��������ȟڟ������$TX_SCREEN 1$�����}��Q�c�u�������?���>�����!� 3�E���ί{������� ÿտL���p��/�A� S�e�w��Ͽ��� �����ߐϢ�O�a� s߅ߗߩ� ���D��� ��'�9�K���o��� ����������d�v� #�5�G�Y�k�}���� ������������C�$UALRM_MSG ?-��:� ;�u� ���� �#�)ZM~q�VS�EV  d��TECFG �&-�7�  ��@�  A! �  B��
  ��-�7/I/[/m// �/�/�/�/�/�/�'��GRP 2'�; 0�	 !/C?�V I_BBL_N�OTE (�T��l��2���V2DEF�PRO` %d (%��?��?�?�? O�?,OOPO;OaO�O�qO�O�O�OL<FKE�YDATA 1)<-�-0p ��0?3_E__i_{_RZ�,(�_�_�([ INST ]�_��^  IRECT �_�_ND�Roo CHOICE�_�;o[EDCMD�Uo�o�PORE�PFO�o�o�o�o�o�o ,>%bI������ ���/frh/gu�i/whitehome.png�`1�C�U�g�y��
�inst�����Џ��􏃇  �direc����9�K�]�o����in������џ������clos���?�Q�c�u������
�edcmd ��.�¯ԯ���
���}
�arwrg�� A�S�e�w�������� ʿܿ� �ϡ�6�H� Z�l�~ϐ�ϴ����� ����ߝ�2�D�V�h� zߌߞ�-��������� 
���@�R�d�v�� ��)���������� *��/�V�h�z����� ����������
. ��Rdv���; ���*<� `r����I� �//&/8/�J/n/ �/�/�/�/�/W/�/�/ ?"?4?F?�/j?|?�? �?�?�?S?�?�?OO 0OBOTO�?xO�O�O�O �O�OaO�O__,_>_ P_�Ob_�_�_�_�_�_ �_o_oo(o:oLo^o��{kk������o�o�m�o�o�o�f,��A( ew^����� ���+��O�6�s� ��l�����͏���� �'��K�]�<����� ����ɟ۟�_���#� 5�G�Y�k��������� ůׯ�x���1�C� U�g�����������ӿ ������-�?�Q�c� u�ϙϫϽ������� ���)�;�M�_�q߃� ߧ߹��������� %�7�I�[�m���� �������������3� E�W�i�{�������� ��������/AS ew��r���� � =Oas ���8���/ /'/�K/]/o/�/�/ �/4/�/�/�/�/?#? 5?�/Y?k?}?�?�?�? B?�?�?�?OO1O�? UOgOyO�O�O�O�OPO �O�O	__-_?_�Oc_ u_�_�_�_�_L_�_�_ oo)o;oMo�_qo�o �o�o�o�oZo�o %7I�om��е��� �{�>� ����� (� �J�\�6�,H��� @�����Տ�Ώ�� /�A�(�e�L������� �������ܟ� �=� $�a�s�Z���~���ͯ ����'�9�K�Z o���������ɿۿj� ���#�5�G�Y��}� �ϡϳ�����f���� �1�C�U�g��ϋߝ� ��������t�	��-� ?�Q�c��߇���� ��������)�;�M� _�q� ����������� ��~�%7I[m ������ �!3EWi{
 ������/� //A/S/e/w/�/��/ �/�/�/�/??�/=? O?a?s?�?�?&?�?�? �?�?OO�?9OKO]O oO�O�O�O4O�O�O�O �O_#_�OG_Y_k_}_ �_�_0_�_�_�_�_o o1o�_Uogoyo�o�o �o>o�o�o�o	- �oQcu���� L����)�;�� _�q���������H�ݏ����%�7�I�  �K��  ���t�����p���̟��,������!��E�W� >�{�b�������կ�� ����/��S�e�L� ��p�����ѿ�ʿ� �+�=�/a�sυϗ� �ϻ�ʏ������'� 9�K���o߁ߓߥ߷� ��X������#�5�G� ��k�}�������� f�����1�C�U��� y�����������b��� 	-?Qc��� �����p );M_���� ����~/%/7/ I/[/m/��/�/�/�/ �/�/z/?!?3?E?W? i?{?Rϟ?�?�?�?�? �? ?O/OAOSOeOwO �OO�O�O�O�O�O_ �O+_=_O_a_s_�__ �_�_�_�_�_oo�_ 9oKo]ooo�o�o"o�o �o�o�o�o�o5G Yk}��0�� �����C�U�g� y�����,���ӏ��� 	��-���Q�c�u��� ����:�ϟ���� )���M�_�q�����������0����0��������*�<��,(�m� ϑ� x���ǿ���ҿ�!� �E�,�i�{�bϟφ� ���ϼ�������A� S�:�w�^ߛ߭ߌ?�� ������+�:�O�a� s�����J����� ��'�9���]�o��� ������F������� #5G��k}�� ��T��1 C�gy���� �b�	//-/?/Q/ �u/�/�/�/�/�/^/ �/??)?;?M?_?�/ �?�?�?�?�?�?l?O O%O7OIO[O�?O�O �O�O�O�O�O��_!_ 3_E_W_i_pO�_�_�_ �_�_�_�_�_o/oAo Soeowoo�o�o�o�o �o�o�o+=Oa s������ ��'�9�K�]�o��� �����ɏۏ���� ��5�G�Y�k�}���� ��şן������1� C�U�g�y�����,��� ӯ���	����?�Q� c�u�����(���Ͽῠ���)� P+�}� P���T�@f�x�PϚϬφ�,�� �ϐ����%�7��[� B�ߑ�xߵߜ����� �����3�E�,�i�P� ��t���������� ��OA�S�e�w����� ����������+ ��Oas���8 ���'�K ]o����F� ��/#/5/�Y/k/ }/�/�/�/B/�/�/�/ ??1?C?�/g?y?�? �?�?�?P?�?�?	OO -O?O�?cOuO�O�O�O �O�O^O�O__)_;_ M_�Oq_�_�_�_�_�_ Z_�_oo%o7oIo[o 2�o�o�o�o�o�o�_ �o!3EWi�o ������v� �/�A�S�e������ ����я������+� =�O�a�s�������� ͟ߟ񟀟�'�9�K� ]�o��������ɯۯ �����#�5�G�Y�k� }������ſ׿��� Ϝ�1�C�U�g�yϋ� ϯ���������	ߘ� -�?�Q�c�u߇ߙ�p`����p`�����������
����,�M� �q�X�� �����������%� �I�[�B��f����� ����������!3 W>{�lo��� ���/ASe w��*���� //�=/O/a/s/�/ �/&/�/�/�/�/?? '?�/K?]?o?�?�?�? 4?�?�?�?�?O#O�? GOYOkO}O�O�O�OBO �O�O�O__1_�OU_ g_y_�_�_�_>_�_�_ �_	oo-o?o�_couo �o�o�o�oLo�o�o );�o_q�� �������%� 7�I�Pm�������� Ǐُh����!�3�E� W��{�������ß՟ d�����/�A�S�e� ����������ѯ�r� ��+�=�O�a�𯅿 ������Ϳ߿񿀿� '�9�K�]�o����ϥ� ��������|��#�5� G�Y�k�}�ߡ߳��� �����ߊ��1�C�U� g�y����������h��	��p���p���4�F�X�0�z���f�,x��p ������;"_ qX�|���� �%I0mT �������� !/3/E/W/i/{/��/ �/�/�/�/�/?�//? A?S?e?w?�??�?�? �?�?�?O�?+O=OOO aOsO�O�O&O�O�O�O �O__�O9_K_]_o_ �_�_"_�_�_�_�_�_ o#o�_GoYoko}o�o �o0o�o�o�o�o �oCUgy��� >���	��-�� Q�c�u�������:�Ϗ ����)�;�/_� q�����������ݟ� ��%�7�I�؟m�� ������ǯV����� !�3�E�ԯi�{����� ��ÿտd�����/� A�S��wωϛϭϿ� ��`�����+�=�O� a��υߗߩ߻����� n���'�9�K�]��� �����������|� �#�5�G�Y�k���� ����������x�@1CUgyP�{��P������������, �-�Q8u�n �����/�)/ ;/"/_/F/�/�/|/�/ �/�/�/??�/7?? [?m?L��?�?�?�?�? �?��O!O3OEOWOiO {O
O�O�O�O�O�O�O �O_/_A_S_e_w__ �_�_�_�_�_�_o�_ +o=oOoaoso�oo�o �o�o�o�o�o'9 K]o��"�� �����5�G�Y� k�}������ŏ׏� ������C�U�g�y� ����,���ӟ���	� ���?�Q�c�u����� ���?ϯ����)� 0�M�_�q��������� H�ݿ���%�7�ƿ [�m�ϑϣϵ�D��� �����!�3�E���i� {ߍߟ߱���R����� ��/�A���e�w�� ������`����� +�=�O���s������� ����\���'9 K]������� �j�#5GY �}��������$UI_INU�SER  ����
!��  ��_M�ENHIST 1�*
%  �(  (/�SOFTPART�/GENLINK�?current�=menupage,153,1)/0�/�/�/�/�)c/u/631�/?1?C?U?' �'�/�.7?�?��?�?�?t6k?�%e�dit�"MAIN�_MANIPULACION�?4OFOXOr�_O�O�O�O�O �O�OmO__&_8_J_ \_�O�_�_�_�_�_�_ i_�_o"o4oFoXojot��Q^!�_�o�o�o �o�o�o�_+=O as����� ���'�9�K�]�o� �������ɏۏ��� ��#�5�G�Y�k�}�� ���şן������ 1�C�U�g�y���vo�o ��ӯ���	���?� Q�c�u�����(���Ͽ ����)ϸ�M�_� qσϕϧ�6������� ��%ߴ�I�[�m�� �ߣߵ�D�������� !�3���W�i�{��� ���������/� A�D�e�w��������� N�����+=O ��s�����\ �'9K�o ������j� /#/5/G/Y/�}/�/ �/�/�/�/����?? 1?C?U?g?j/�?�?�? �?�?�?t?�?O-O?O QOcOuOO�O�O�O�O �O�O�O_)_;_M___ q_ __�_�_�_�_�_ o�_%o7oIo[omoo o�o�o�o�o�o�o�/���$UI_PA�NEDATA 1�,���3q�  	�}�/frh/gu�iJqdev0.s�tm ?_wid�th=0&_height=10cp�Rpice=TP&�_lines=1�5&_colum�ns=4cpfon�t=24&_pa�ge=whole�Rp�&)pri9m��  }��`�&�8�J�\� )^� ��i�����ʏ܏Ï � �$�6��Z�A�~����w����&�� �    I�����'� 9�K���o�������� ɯۯ�T��#�
�G� .�k�}�d�����ſ׿ ������1��U�ȗ 6pt�5s���ϧϹ� ������B�߆�7�I� [�m�ߑ��ϵ��߮� �����!��E�,�i� P����������� l�~�/�A�S�e�w��� ��� ������� +=��aH�l� �����9  ]oV���� ���/#/vG/Y/ ��}/�/�/�/�/�/>/ �/�/?1??U?<?y? �?r?�?�?�?�?�?	O �?-O��p/uO�O�O �O�O�O"O�Of/_)_ ;_M___q_�O�_�_�_ �_�_�_o�_%ooIo 0omoofo�o�o�o�o LO^O!3EWi �o� _����� ���A�(�e�L��� �����������܏�  �=�O�6�s��o�o�� ��͟ߟ��V�'�9� �]�o���������� ۯ¯�����5��Y� k�R���v���ſ���0пπ���}��W� i�{ύϟϱ�)E��� I�����&�8�J�\� �π�gߤߋߝ����� ����"�4��X�?�|����u��B������$�UI_POSTY�PE  ��� 	 ������QUICKM_EN  �������RESTOR�E 1-��  ���BK������K�m�� ����+��Oa s��:���� ��"4�o� ���Z���/ #/5/�Y/k/}/�/�/ L�/�/�/D/??1? C?U?�/y?�?�?�?�? d?�?�?	OO-O�/�? LO^O�?�O�O�O�O�O �O�O_)_;_M____ �_�_�_�_�_vO�_�_ �_n_7oIo[omoo"o �o�o�o�o�o�o�o!�3EWi#�SCR�E3�?8��u1sc��u2��t3�t4�t5�t6ʤt7�t8�q�sTAT��� G���USER�p��rTL�p�sks�s?�4?�U5?�6?�7?�8?����NDO_CFG� .��.�-���P�D�q!��?None ����_INFO 1/j��ˀE�0%o �B�ԏ���9�K�.� o���d�����ɟ۟��������5����OFFSET 2��ρB�
s}����� ���������(� r�,�y�p��������� �ܿ� �J�H�L�:��o�
_ϔ�N�UFR�AME  
t�����RTOL_A�BRT��R���EN�B����GRP 1�3x�D�Cz  A�/�-э�-�?�Q߀c�u߇ߙ߫���2�U��ȍ���MSK  ���ˁ��N��%�É�%�=�%�VC�MR�29d����p	�� ��1: SC130EF2 *���
te�I�����Ԃ5p���?���@��p:���A� ������x�,�Y�~�T��������A�r�m���r B�����q��e���E� "��F1jU�y ������0���TfO�ISIO�NTMOU����懅�}y�:SﳸS� $� FR:\�\��A\k �߀ MC�LO�G�   UD�1�EX�q'� B@ �� 2"!,�P/!T/x/
s� � n6  ���v/"����`�&�  =����!
t�  }�TRAIN/��"�"��  d
3Qp�)�Z�;d�( �%J=J?X?j?|?�? �?�?�?�?�?�?OOh0OBOw_ RE��<ل�O�LEXEr�=d���1-em�VMPHAS�p䠅����P�RTD�_FILTER �2>d� �L�� ��5_G_Y_k_}_�_�_ �_�_�_G�#_oo,o >oPoboto�o�o�oM��SHIFT��1?d�
 <?,+� �u�o	B+xO a��������,���b�9�	L�IVE/SNAP��vsfliv\�Nt�� ^�yU����menu�����L��#����e�@X�i	�eMO�A�N�ĺ��$WAIT?DINEND��؂��O���ߡ����S�˟��TIM������G�����;�ʟ�������REL�E�A�π�����_ACT��ʨ���� B�%�K������RDIS���ρ�V�_AXSR��2C��]�^�V*1_IoR  J� �� ѿ�����+�=�O� a�sυϗϩϻ����� ����'�9�K�]�o� �ߓߥ߷��������� �#�5�G�Y�k�}���������|XVR�f�D�N�$ZA�BC*21E�K �,0 2��oZI-P�F�O�������G�MPCF_/G 1G��04q�������H���S ��E@<�P Ju6�Z?�7������4�gyG �=���� ������@I]��U�YLINDQJ �> ,(  *O/`-EL/0�/p/�/�- b�/ �/>I/*?�/N?5?G? �?�/�?�?�??�?�? q?&OOJO1O�?�O�O�F�2K��� ����O�Lʳa__�:_>�Oj_>��QA��$SPHERE 2L/-��?�_4O �_�_�_obOu_Pobo �?�o%oo�o�o�o�o 9o(oo�o^�o� i{��o�� ��ZZ� �R�