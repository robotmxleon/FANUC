��   m�A��*SYST�EM*��V9.0�055 1/3�1/2017 �A   ����DMR_GRP�_T  � �$MA��R_D�ONE  $�OT_MINUS�   	GPyLN8COUNP �T REF>wP�OOtlTpB�CKLSH_SI�GoSEACHMsST>pSPC�
��MOVB RAD�APT_INERzP �FRIC�
_COL_P M�
�GRAV��� HsIS��DSP?��HIFT_ER[RO�  �NA�pMCHY SwARM_PARA#w d7ANGC �M2pCLDE|�CALIB� �DB$GEARz�2� RING���<$1_8k/�<�FMS*�t *v M_LIF��u,(8*���M(DSTB0+_0>*_���*#z&~+CL_TIM��PCCOMi�F�Bk M� �MAL�_�EC�S�P�!Q%XO g$PS� �TI����%�"r $DT�Y?R. l*1EN�D14�$1�ACT�1#4V22\93\94�\95\96\6_OVR\6� GA[7�2h7 �2u7�2�7�2�7�2�8oFRMZ\6DE�{DX\6CURL� 
HSZ27Fh1DGu1�DG�1DG�1DG�1DCN�A!1?( �P�L� + ��S�TA23TRQ_Mȫ�/@K"�FSX��JY�JZ�II�JI��JI�D �$U1S�S  ����6Q����+PVE�RSI� 4W�  ��GQIRTUAL3_EQ'� 1 TX + ��(P���_ �_�_�_o�_%oo"o�[oFoojjAQ�o�l�������K����/ 舡�[������o �o�o�l/VSe�k��r�������d�#�5�G����=L��R�y�?�z���@�����я �����+�=�O�a�s���� rU����8��ޟ:T  2�� !�3�E�W�i�{���������<��ۯ���� #�5�G�Y�k�}��������sP��$$ 1��\�qF�6 F@���� 
Ϙ��@�+�d�Oψ� sϬϗϼ�������π*��N�9�K߄��� ��ߓ�t������� r�7���[�m��>�P� ����������!�3� ��W�i�{�:�L����� ������/��S ew6H���� �+�Oas 2D�����/ /'/�K/]/o/./@/ �/�/�/�/�/�/?�� ;Q�/K?]?o?�/�?�? �?�?�?�?�?O#O�? GOYOkO*O�O�O�O�O �O�O�O__�OC_U_�g_��,($1234567890�_ �U���_�_�_�_�_�_ oo;o+oGoOoao�o �o�o�o�o�o�o�o I9U]y�� �����!��-� 5�G�{�k�������Տ~Ņ�$PLCLų��� �D!�?�   �1�%�T�!�x�c��� ������������� >�P�