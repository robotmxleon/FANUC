��   F��A��*SYST�EM*��V9.0�055 1/3�1/2017 ?A #  �����#�AMON_D�O_T   �$PORT_�TYPE  �@NUMJ/SG�NL7 L�$MIN_RAN}GI$MAXr�NOo ALxp V��~ �COUNT>J��AWE08 �� $AWn0ENBJ $�|G1LY_TIV�$WRN_ALM�STP�
�E��C�.�WT�C�
J�AFT_�CHGxAVRG�_INT��{SgAVE�YP1?ER_REG�Tw$WA� SIG�� OP��V/OLTS�����AMP�&AEx �#E_VL� �&D'>% I*f$� _�ANL�  �p 
$US0 S�_CMD � PRIORITY�"�UPPER� $�LOW�$�#$FgDBK�"�RAv ~�!SQ_AVG�#n�#SD_� CE� 8� ��$ �� � �LIN�!$ARC_ENABL�!|� 0DETEC�!~< ELD_SP�$?PD_UNI��!N92DIS�"�ID sIM�#�� l v1WFt2θ�CF�" � �$PS_MANU�F �2OD�EL�5PROCEySN0�0WFEEW0�ESC�2�2_FI�#1�1�1�7T _AOT�"�2I�6D�7DC`1�6L �"{2 � �CNV� 7   $EQ�zx�ODOU��2?@T�Bd  $~?C 2 kE�DD   , �� MM�!�$D� ��!2� $F� �B�4NuV7	JBSEL10�_NOJDATA�_s@�@ �2W�PpG
{M
�FWP�7 L@�L
 ��WIR_CLP4 L@AS�BU8  H $(4��R�4��YPREF� �U �}!ECU��  �JB~ �S  � $BPEEPf#�}!SCH7 � �!��`�1e�#dPK*jFRE�Q.gULSwbSP�0fg2y�!hyb�*g�F�"AI6 �ZCoVG}�hp dD��e�e�`�	�a��dBzVB�aZEROy�}uSLO]R�`NT�!P�cO	U\93��L FORMA0NqAra�0J3	� �D�cQWUXWE�IOEX74� �A�Wfxcc�pS_91INp�� :1�U�p� FAU�G"t0LO�0�qPD�!�G��R<�ADp�;�STIC�@�pR�OBOT�ADY��rERRO�SE���`S��p�!TR���$S�CHDOG�_�@%��0_ACTSIV���I�C�0�1�2�q�OTF~7 � $
� �P��x�nfpNCi0�c;�f0� *d;�*g0�7f;�7i0��Fd;�Fg~�Td��TfU�P�@�B:BEPCR�7�� WSTK��� =�Hr ՒƁ %��00��2�X���0�A~�3KIPTH�E91�S;������PIKEf���0�0�WWV�2t�E_HaO;0�0��PHK-18���� RMT����SPTL�0p�$�Hz��SW��pd�$BBg1_ONL4�$B�2pf�bgF�WF�1e2_R��0zE"�!� _W;6�A?ND1OFF���!�ND2g�3g�R�Sp� �A� jCEPM�? | $�0�@ g��e��*f��7b���Ff�TfADAPTz� G�CSENS��c��!ݒ��8 � 0?,2���"��$ �1b�!c�7cc�Fa|� Tac�^��'y��&l��&*�!4�&5�&6�"8��W�@�2 HOU�!h�o � �SE�0 �g4�Q�T<��6��'��46�q56�0� ?%$CURR7(�^�"HEATzPe@ �!燰"j���i�p��GAP�#Ti�XPY0���EHP��@��pDS��@�!GP�0S�!�$���$GO� RI����AM�#/"�#M䩰jAN3O�BEFB ;�LHV1[5j�� 43;1 `H�V�PA�H�r���3��F1�� �D�POSR 7 W� 	� RSB�$ ��0G�m�b�O�J���,O��DU�IW�AXQl�2C,1L�"!D����?3|!E��8  4�@P֋q]��SGʦ�~�;A8�8 ? $ $�@�CL�$��s	�R|��$ ;o2� �"��ql��q��� 	PK �P��
��*���q@�Ba��b�@4�5�6:2K�3������FW�q�B<��ALAR���2 ��2�����
�3�Q_R}��
`�.44�F�+�PW,���_@ĸ�Ӕ]� ������Qbwm��t���QDI�c�j��p~pus�R�SIZ���BOAR���1]E7�]�\�h"�0h"��ķ�$V�END��I��DE'VIC��0D�����MAJ��V�#IN`�(�$�uI"�vMA���pFI�0�BW��b�E�� p $@��X�� ⡡��F̀OR_R��C�^1D4gTO_��O5_R�p3RS<�'�OS�9�r�UP� # N�:��0�`�=� �6�x�6��9PURG�,�RKtSTFR�p&���A��.E�.E� AED��P-��M%�fM!T�����eEM7��Q �5���Z$�22�9�P�駇��K�p�QADJ��T��NEXT��r_LE�c��P��X��AM����aA��_�#�IV���H�q�2�eFL������P��:���`�0�8� ��;�WT[�6��CY�� ��  �	`��`�( �bTOTAL_��Q�c���VI�p�WW#ARo��U��A*�bPY&1b�uKG����'" A}�#N�p � �aSCFG�1z�LOO�B:��P�Q�S!@�<��GLOB�P�⸣�� ��NOT���$0QI4�*��AVh�Y��$�������|�e��W_SHFL�%W�X�fkrI�$�q �e�RY	��оP8��%�ʀLIMS`�i��@�c7�UIF�e�APCOUPL�R @ �p�q���� �qUR�`N:��<�MMYm �u�0�u�  ����U�STOk�   � x�0 �qp`� 
  ��SEM�Gg��1! ,��M�G�Ag���NOzPR� ����wa�"� ,/���Ȣ=6Ƞ��3T� )�RT���p�`��=����AHER� ��A�������'"݈{ �������@���Q�L� �)BD ��2C���7B�<�i3_FIL@�Wn��BUG_3SM ���ñF_F����q�4, _4N SV@БT�C�P��=Ҕ�DIO�������.a�3TM�C��PA�Pq���qw�x��q�_DY�NV�2Wԣ����KEYV�GQׂ���F��?�/B�{�_C:��R�TOU����8�Б��CAL�Q0D�`� TIp1�P_y��RT���@��A?2��$$CLAS�S  ���4���� �-��SB��� � ���IRT�U�����AWAOLY1�� 
��$��
�K���n�2�f�[�[���g�
�?�������g� ����������(π:�L�^�pςϑ�l�EXEu�`��������� Ͽ�*�<�N�`�r߄���ߨߺߕ�r@S Rw���:����#�5� G�Y�k�}���������������l�NLoG 2x� ��ߊ��?��<1�6�`���e��� p`����{` �2:�)��General� Purpose��MIG (Volts, 0�)��� ����
A�WMGENL.V�RA*EGLGMG19��g�` ��������'���� �����������CNV 2	x�=�[����� 4aPzU h�����// �=/O/./s/�/\�/ �/b/�/�/�/?'?? K?]?<?�?�?r?�?�� E�/�?O�?2ODO#O hOzOYO�O�O�O�O�O �O
__�?@_R_�Ov_ �_g_�_�_�_�_�_�_ o�_(oNo�?ro-_�o �o3o�o�o�o�o 8J)nM_�{o ������ �F� %�j�|�[�������֏ �go���0�B�!�f� E�W���{���ҟ���� ��,�>��b�t�� ������ί௿��� ��:�L�+�p����O� ��ʿU�� �߿$�6� �Z�l�KϐϢρ��� �ϯ���ߵ�2�D�#� h�z�Yߞ�}ߏ��߳����
��NVWP �2|	i\>�T �
��b�t���US�TOM 2|l  ���������h�	hd"���DEFSCH R|��Q�<�b�@D�efault Schg���n������� ����K"4 �Xj��������
)�FBKLO_G1 @��T����  Ugy��12=O�����5LG_CNT�  ����)�IO_EX 2�����[A ��C�]$@�������!�
W�eld Spee�%��IPM   d$�/�/�/�/??(?�:?��OTF 2��A?�?�?�?�?��?C8=�����@᠛��?K)�PCR� 2��pI�BH�?��BC!�FK<D7��*����?�ffAAZ �A"��OFM"@����/�O@uO"@����9�WOELG��k%*_��F�023456�78901JRUK% 4_y_�_�_HIȩ_7]��OOSRAM2���IB�$�_oCRG�SEL R<��Q� 	Process 1oSf�2�_oj3i�o4
i�o5�-mlXS���o7��kn8i�'l"@��� 1�_);Es-B� �W��%VoltWage��qsf�c%Dw|!@]�y�h��aW�ire f�  s�$	� hc%[&t/ �oDS�l*�<�N�`� r���������̏ޏ��@��&�]+zvd"�����  �#��E�Z"!��a��^/�� ��V���a�a�ɒCurre{nt�Amp� =���l�eu���Q�c� u���������ϯ�� ��)�;�M��W���a �����ឱ	q��)q�� Iq��R�͹ϧg�a�a A��b-���-�	q-�)qH-�VE!��\e�	q_?���*�Z�% ������ϻ�����ߜPDRuS R\zH�A�jq��C�U�g��� ��gߩ߻�u߇ߙ�� �������]�o�)�;� M��������#� �����k�}�7�I�[� ����������1C ��I��Wi� �����?Q /������ //)/;/M+�U/g) {/�/�/M/�/?cS2�S�^=R��b�S2U�PYp^=�=�_o?�33H1>E0�=L��>I0h!*�@"�@#�@$�1t9&�g�q�#?�v�#�>�8�8CWIRE 2&M<�?�?h��>�3�>�G�(=�J*�ESCFG �G�A���Y��OOˎE7])COWUPL�0=k
0�vkB`�D�^�L�[ �OZW�O�G_�OP_G_|Y\�HNB  ���Ec&FUSTOM  =k
8ƙy�O&E�EMGOFF �!=kS��)BPC�R "�_��@���zqC{sUūMJo�\ zt�f_oeo��
Cl� q¨1